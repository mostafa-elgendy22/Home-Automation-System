/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Mon Dec 20 17:51:29 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1771793495 */

module first_stage(A, B, clk, enable, negative_product_second_stage, 
      next_stage_enable, operand1, operand2);
   input [15:0]A;
   input [15:0]B;
   input clk;
   input enable;
   output negative_product_second_stage;
   output next_stage_enable;
   output [14:0]operand1;
   output [14:0]operand2;

   wire n_0_0;
   wire n_0_29;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_14;
   wire n_0_0_3;
   wire n_0_15;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_16;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_17;
   wire n_0_0_8;
   wire n_0_18;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_19;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_20;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_21;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_22;
   wire n_0_0_17;
   wire n_0_23;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_24;
   wire n_0_0_20;
   wire n_0_25;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_26;
   wire n_0_0_23;
   wire n_0_27;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_1;
   wire n_0_0_27;
   wire n_0_2;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_3;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_4;
   wire n_0_0_32;
   wire n_0_5;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_6;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_7;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_8;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_9;
   wire n_0_0_41;
   wire n_0_10;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_11;
   wire n_0_0_44;
   wire n_0_12;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_13;
   wire n_0_0_47;
   wire n_0_28;

   DFF_X1 \operand2_reg[14]  (.D(n_0_28), .CK(n_0_0), .Q(operand2[14]), .QN());
   DFF_X1 \operand2_reg[13]  (.D(n_0_13), .CK(n_0_0), .Q(operand2[13]), .QN());
   DFF_X1 \operand2_reg[12]  (.D(n_0_12), .CK(n_0_0), .Q(operand2[12]), .QN());
   DFF_X1 \operand2_reg[11]  (.D(n_0_11), .CK(n_0_0), .Q(operand2[11]), .QN());
   DFF_X1 \operand2_reg[10]  (.D(n_0_10), .CK(n_0_0), .Q(operand2[10]), .QN());
   DFF_X1 \operand2_reg[9]  (.D(n_0_9), .CK(n_0_0), .Q(operand2[9]), .QN());
   DFF_X1 \operand2_reg[8]  (.D(n_0_8), .CK(n_0_0), .Q(operand2[8]), .QN());
   DFF_X1 \operand2_reg[7]  (.D(n_0_7), .CK(n_0_0), .Q(operand2[7]), .QN());
   DFF_X1 \operand2_reg[6]  (.D(n_0_6), .CK(n_0_0), .Q(operand2[6]), .QN());
   DFF_X1 \operand2_reg[5]  (.D(n_0_5), .CK(n_0_0), .Q(operand2[5]), .QN());
   DFF_X1 \operand2_reg[4]  (.D(n_0_4), .CK(n_0_0), .Q(operand2[4]), .QN());
   DFF_X1 \operand2_reg[3]  (.D(n_0_3), .CK(n_0_0), .Q(operand2[3]), .QN());
   DFF_X1 \operand2_reg[2]  (.D(n_0_2), .CK(n_0_0), .Q(operand2[2]), .QN());
   DFF_X1 \operand2_reg[1]  (.D(n_0_1), .CK(n_0_0), .Q(operand2[1]), .QN());
   DFF_X1 \operand2_reg[0]  (.D(B[0]), .CK(n_0_0), .Q(operand2[0]), .QN());
   DFF_X1 \operand1_reg[14]  (.D(n_0_27), .CK(n_0_0), .Q(operand1[14]), .QN());
   DFF_X1 \operand1_reg[13]  (.D(n_0_26), .CK(n_0_0), .Q(operand1[13]), .QN());
   DFF_X1 \operand1_reg[12]  (.D(n_0_25), .CK(n_0_0), .Q(operand1[12]), .QN());
   DFF_X1 \operand1_reg[11]  (.D(n_0_24), .CK(n_0_0), .Q(operand1[11]), .QN());
   DFF_X1 \operand1_reg[10]  (.D(n_0_23), .CK(n_0_0), .Q(operand1[10]), .QN());
   DFF_X1 \operand1_reg[9]  (.D(n_0_22), .CK(n_0_0), .Q(operand1[9]), .QN());
   DFF_X1 \operand1_reg[8]  (.D(n_0_21), .CK(n_0_0), .Q(operand1[8]), .QN());
   DFF_X1 \operand1_reg[7]  (.D(n_0_20), .CK(n_0_0), .Q(operand1[7]), .QN());
   DFF_X1 \operand1_reg[6]  (.D(n_0_19), .CK(n_0_0), .Q(operand1[6]), .QN());
   DFF_X1 \operand1_reg[5]  (.D(n_0_18), .CK(n_0_0), .Q(operand1[5]), .QN());
   DFF_X1 \operand1_reg[4]  (.D(n_0_17), .CK(n_0_0), .Q(operand1[4]), .QN());
   DFF_X1 \operand1_reg[3]  (.D(n_0_16), .CK(n_0_0), .Q(operand1[3]), .QN());
   DFF_X1 \operand1_reg[2]  (.D(n_0_15), .CK(n_0_0), .Q(operand1[2]), .QN());
   DFF_X1 \operand1_reg[1]  (.D(n_0_14), .CK(n_0_0), .Q(operand1[1]), .QN());
   DFF_X1 \operand1_reg[0]  (.D(A[0]), .CK(n_0_0), .Q(operand1[0]), .QN());
   DFF_X1 negative_product_second_stage_reg (.D(n_0_29), .CK(n_0_0), .Q(
      negative_product_second_stage), .QN());
   CLKGATETST_X1 clk_gate_operand2_reg (.CK(clk), .E(enable), .SE(1'b0), 
      .GCK(n_0_0));
   XOR2_X1 i_0_0_0 (.A(A[15]), .B(B[15]), .Z(n_0_29));
   NAND2_X1 i_0_0_1 (.A1(A[15]), .A2(enable), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_0), .ZN(n_0_0_1));
   NAND2_X1 i_0_0_3 (.A1(n_0_0_1), .A2(A[0]), .ZN(n_0_0_2));
   XNOR2_X1 i_0_0_4 (.A(n_0_0_2), .B(A[1]), .ZN(n_0_14));
   OAI21_X1 i_0_0_5 (.A(n_0_0_1), .B1(A[1]), .B2(A[0]), .ZN(n_0_0_3));
   XNOR2_X1 i_0_0_6 (.A(n_0_0_3), .B(A[2]), .ZN(n_0_15));
   INV_X1 i_0_0_7 (.A(n_0_0_3), .ZN(n_0_0_4));
   AOI21_X1 i_0_0_8 (.A(n_0_0_4), .B1(A[2]), .B2(n_0_0_1), .ZN(n_0_0_5));
   XNOR2_X1 i_0_0_9 (.A(n_0_0_5), .B(A[3]), .ZN(n_0_16));
   OAI21_X1 i_0_0_10 (.A(n_0_0_1), .B1(A[3]), .B2(A[2]), .ZN(n_0_0_6));
   NAND2_X1 i_0_0_11 (.A1(n_0_0_3), .A2(n_0_0_6), .ZN(n_0_0_7));
   XOR2_X1 i_0_0_12 (.A(n_0_0_7), .B(A[4]), .Z(n_0_17));
   AOI21_X1 i_0_0_13 (.A(n_0_0_7), .B1(A[4]), .B2(n_0_0_1), .ZN(n_0_0_8));
   XNOR2_X1 i_0_0_14 (.A(n_0_0_8), .B(A[5]), .ZN(n_0_18));
   INV_X1 i_0_0_15 (.A(n_0_0_8), .ZN(n_0_0_9));
   AOI21_X1 i_0_0_16 (.A(n_0_0_9), .B1(A[5]), .B2(n_0_0_1), .ZN(n_0_0_10));
   XNOR2_X1 i_0_0_17 (.A(n_0_0_10), .B(A[6]), .ZN(n_0_19));
   INV_X1 i_0_0_18 (.A(n_0_0_10), .ZN(n_0_0_11));
   AOI21_X1 i_0_0_19 (.A(n_0_0_11), .B1(A[6]), .B2(n_0_0_1), .ZN(n_0_0_12));
   XNOR2_X1 i_0_0_20 (.A(n_0_0_12), .B(A[7]), .ZN(n_0_20));
   INV_X1 i_0_0_21 (.A(n_0_0_12), .ZN(n_0_0_13));
   AOI21_X1 i_0_0_22 (.A(n_0_0_13), .B1(A[7]), .B2(n_0_0_1), .ZN(n_0_0_14));
   XNOR2_X1 i_0_0_23 (.A(n_0_0_14), .B(A[8]), .ZN(n_0_21));
   INV_X1 i_0_0_24 (.A(A[8]), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_25 (.A(n_0_0_14), .B1(n_0_0_15), .B2(n_0_0_0), .ZN(n_0_0_16));
   XOR2_X1 i_0_0_26 (.A(n_0_0_16), .B(A[9]), .Z(n_0_22));
   AOI21_X1 i_0_0_27 (.A(n_0_0_16), .B1(A[9]), .B2(n_0_0_1), .ZN(n_0_0_17));
   XNOR2_X1 i_0_0_28 (.A(n_0_0_17), .B(A[10]), .ZN(n_0_23));
   INV_X1 i_0_0_29 (.A(A[10]), .ZN(n_0_0_18));
   OAI21_X1 i_0_0_30 (.A(n_0_0_17), .B1(n_0_0_18), .B2(n_0_0_0), .ZN(n_0_0_19));
   XOR2_X1 i_0_0_31 (.A(n_0_0_19), .B(A[11]), .Z(n_0_24));
   AOI21_X1 i_0_0_32 (.A(n_0_0_19), .B1(A[11]), .B2(n_0_0_1), .ZN(n_0_0_20));
   XNOR2_X1 i_0_0_33 (.A(n_0_0_20), .B(A[12]), .ZN(n_0_25));
   INV_X1 i_0_0_34 (.A(A[12]), .ZN(n_0_0_21));
   OAI21_X1 i_0_0_35 (.A(n_0_0_20), .B1(n_0_0_21), .B2(n_0_0_0), .ZN(n_0_0_22));
   XOR2_X1 i_0_0_36 (.A(n_0_0_22), .B(A[13]), .Z(n_0_26));
   AOI21_X1 i_0_0_37 (.A(n_0_0_22), .B1(A[13]), .B2(n_0_0_1), .ZN(n_0_0_23));
   XNOR2_X1 i_0_0_38 (.A(n_0_0_23), .B(A[14]), .ZN(n_0_27));
   NAND2_X1 i_0_0_39 (.A1(B[15]), .A2(enable), .ZN(n_0_0_24));
   INV_X1 i_0_0_40 (.A(n_0_0_24), .ZN(n_0_0_25));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_25), .A2(B[0]), .ZN(n_0_0_26));
   XNOR2_X1 i_0_0_42 (.A(n_0_0_26), .B(B[1]), .ZN(n_0_1));
   OAI21_X1 i_0_0_43 (.A(n_0_0_25), .B1(B[1]), .B2(B[0]), .ZN(n_0_0_27));
   XNOR2_X1 i_0_0_44 (.A(n_0_0_27), .B(B[2]), .ZN(n_0_2));
   INV_X1 i_0_0_45 (.A(n_0_0_27), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_46 (.A(n_0_0_28), .B1(B[2]), .B2(n_0_0_25), .ZN(n_0_0_29));
   XNOR2_X1 i_0_0_47 (.A(n_0_0_29), .B(B[3]), .ZN(n_0_3));
   OAI21_X1 i_0_0_48 (.A(n_0_0_25), .B1(B[3]), .B2(B[2]), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_49 (.A1(n_0_0_27), .A2(n_0_0_30), .ZN(n_0_0_31));
   XOR2_X1 i_0_0_50 (.A(n_0_0_31), .B(B[4]), .Z(n_0_4));
   AOI21_X1 i_0_0_51 (.A(n_0_0_31), .B1(B[4]), .B2(n_0_0_25), .ZN(n_0_0_32));
   XNOR2_X1 i_0_0_52 (.A(n_0_0_32), .B(B[5]), .ZN(n_0_5));
   INV_X1 i_0_0_53 (.A(n_0_0_32), .ZN(n_0_0_33));
   AOI21_X1 i_0_0_54 (.A(n_0_0_33), .B1(B[5]), .B2(n_0_0_25), .ZN(n_0_0_34));
   XNOR2_X1 i_0_0_55 (.A(n_0_0_34), .B(B[6]), .ZN(n_0_6));
   INV_X1 i_0_0_56 (.A(n_0_0_34), .ZN(n_0_0_35));
   AOI21_X1 i_0_0_57 (.A(n_0_0_35), .B1(B[6]), .B2(n_0_0_25), .ZN(n_0_0_36));
   XNOR2_X1 i_0_0_58 (.A(n_0_0_36), .B(B[7]), .ZN(n_0_7));
   INV_X1 i_0_0_59 (.A(n_0_0_36), .ZN(n_0_0_37));
   AOI21_X1 i_0_0_60 (.A(n_0_0_37), .B1(B[7]), .B2(n_0_0_25), .ZN(n_0_0_38));
   XNOR2_X1 i_0_0_61 (.A(n_0_0_38), .B(B[8]), .ZN(n_0_8));
   INV_X1 i_0_0_62 (.A(B[8]), .ZN(n_0_0_39));
   OAI21_X1 i_0_0_63 (.A(n_0_0_38), .B1(n_0_0_39), .B2(n_0_0_24), .ZN(n_0_0_40));
   XOR2_X1 i_0_0_64 (.A(n_0_0_40), .B(B[9]), .Z(n_0_9));
   AOI21_X1 i_0_0_65 (.A(n_0_0_40), .B1(B[9]), .B2(n_0_0_25), .ZN(n_0_0_41));
   XNOR2_X1 i_0_0_66 (.A(n_0_0_41), .B(B[10]), .ZN(n_0_10));
   INV_X1 i_0_0_67 (.A(B[10]), .ZN(n_0_0_42));
   OAI21_X1 i_0_0_68 (.A(n_0_0_41), .B1(n_0_0_42), .B2(n_0_0_24), .ZN(n_0_0_43));
   XOR2_X1 i_0_0_69 (.A(n_0_0_43), .B(B[11]), .Z(n_0_11));
   AOI21_X1 i_0_0_70 (.A(n_0_0_43), .B1(B[11]), .B2(n_0_0_25), .ZN(n_0_0_44));
   XNOR2_X1 i_0_0_71 (.A(n_0_0_44), .B(B[12]), .ZN(n_0_12));
   INV_X1 i_0_0_72 (.A(B[12]), .ZN(n_0_0_45));
   OAI21_X1 i_0_0_73 (.A(n_0_0_44), .B1(n_0_0_45), .B2(n_0_0_24), .ZN(n_0_0_46));
   XOR2_X1 i_0_0_74 (.A(n_0_0_46), .B(B[13]), .Z(n_0_13));
   AOI21_X1 i_0_0_75 (.A(n_0_0_46), .B1(B[13]), .B2(n_0_0_25), .ZN(n_0_0_47));
   XNOR2_X1 i_0_0_76 (.A(n_0_0_47), .B(B[14]), .ZN(n_0_28));
endmodule

module datapath__0_4(operand2, operand1, mult);
   input [14:0]operand2;
   input [14:0]operand1;
   output [29:0]mult;

   HA_X1 i_0 (.A(n_617), .B(n_781), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(n_605), .B(n_616), .CI(n_629), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(n_640), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(n_592), .B(n_604), .CI(n_615), .CO(n_7), .S(n_6));
   FA_X1 i_4 (.A(n_628), .B(n_639), .CI(n_5), .CO(n_9), .S(n_8));
   HA_X1 i_5 (.A(n_3), .B(n_8), .CO(n_11), .S(n_10));
   FA_X1 i_6 (.A(n_579), .B(n_591), .CI(n_603), .CO(n_13), .S(n_12));
   FA_X1 i_7 (.A(n_614), .B(n_627), .CI(n_638), .CO(n_15), .S(n_14));
   FA_X1 i_8 (.A(n_7), .B(n_9), .CI(n_14), .CO(n_17), .S(n_16));
   HA_X1 i_9 (.A(n_12), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_10 (.A(n_567), .B(n_578), .CI(n_590), .CO(n_21), .S(n_20));
   FA_X1 i_11 (.A(n_602), .B(n_613), .CI(n_626), .CO(n_23), .S(n_22));
   FA_X1 i_12 (.A(n_637), .B(n_15), .CI(n_13), .CO(n_25), .S(n_24));
   FA_X1 i_13 (.A(n_22), .B(n_20), .CI(n_24), .CO(n_27), .S(n_26));
   HA_X1 i_14 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_15 (.A(n_553), .B(n_566), .CI(n_577), .CO(n_31), .S(n_30));
   FA_X1 i_16 (.A(n_589), .B(n_601), .CI(n_612), .CO(n_33), .S(n_32));
   FA_X1 i_17 (.A(n_625), .B(n_636), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_18 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_19 (.A(n_32), .B(n_30), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_20 (.A(n_36), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_21 (.A(n_540), .B(n_552), .CI(n_565), .CO(n_43), .S(n_42));
   FA_X1 i_22 (.A(n_576), .B(n_588), .CI(n_600), .CO(n_45), .S(n_44));
   FA_X1 i_23 (.A(n_611), .B(n_624), .CI(n_635), .CO(n_47), .S(n_46));
   FA_X1 i_24 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_48));
   FA_X1 i_25 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_51), .S(n_50));
   FA_X1 i_26 (.A(n_48), .B(n_37), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_27 (.A(n_39), .B(n_50), .CO(n_55), .S(n_54));
   FA_X1 i_28 (.A(n_528), .B(n_539), .CI(n_551), .CO(n_57), .S(n_56));
   FA_X1 i_29 (.A(n_564), .B(n_575), .CI(n_587), .CO(n_59), .S(n_58));
   FA_X1 i_30 (.A(n_599), .B(n_610), .CI(n_623), .CO(n_61), .S(n_60));
   FA_X1 i_31 (.A(n_634), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_32 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_64));
   FA_X1 i_33 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_67), .S(n_66));
   FA_X1 i_34 (.A(n_51), .B(n_64), .CI(n_66), .CO(n_69), .S(n_68));
   HA_X1 i_35 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_36 (.A(n_514), .B(n_527), .CI(n_538), .CO(n_73), .S(n_72));
   FA_X1 i_37 (.A(n_550), .B(n_563), .CI(n_574), .CO(n_75), .S(n_74));
   FA_X1 i_38 (.A(n_586), .B(n_598), .CI(n_609), .CO(n_77), .S(n_76));
   FA_X1 i_39 (.A(n_622), .B(n_633), .CI(n_61), .CO(n_79), .S(n_78));
   FA_X1 i_40 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_81), .S(n_80));
   FA_X1 i_41 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_83), .S(n_82));
   FA_X1 i_42 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_85), .S(n_84));
   FA_X1 i_43 (.A(n_67), .B(n_82), .CI(n_84), .CO(n_87), .S(n_86));
   HA_X1 i_44 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_45 (.A(n_500), .B(n_513), .CI(n_526), .CO(n_91), .S(n_90));
   FA_X1 i_46 (.A(n_537), .B(n_549), .CI(n_562), .CO(n_93), .S(n_92));
   FA_X1 i_47 (.A(n_573), .B(n_585), .CI(n_597), .CO(n_95), .S(n_94));
   FA_X1 i_48 (.A(n_608), .B(n_621), .CI(n_632), .CO(n_97), .S(n_96));
   FA_X1 i_49 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_99), .S(n_98));
   FA_X1 i_50 (.A(n_79), .B(n_96), .CI(n_94), .CO(n_101), .S(n_100));
   FA_X1 i_51 (.A(n_92), .B(n_90), .CI(n_81), .CO(n_103), .S(n_102));
   FA_X1 i_52 (.A(n_98), .B(n_83), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_53 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_54 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   FA_X1 i_55 (.A(n_488), .B(n_499), .CI(n_512), .CO(n_111), .S(n_110));
   FA_X1 i_56 (.A(n_525), .B(n_536), .CI(n_548), .CO(n_113), .S(n_112));
   FA_X1 i_57 (.A(n_561), .B(n_572), .CI(n_584), .CO(n_115), .S(n_114));
   FA_X1 i_58 (.A(n_596), .B(n_607), .CI(n_620), .CO(n_117), .S(n_116));
   FA_X1 i_59 (.A(n_631), .B(n_97), .CI(n_95), .CO(n_119), .S(n_118));
   FA_X1 i_60 (.A(n_93), .B(n_91), .CI(n_99), .CO(n_121), .S(n_120));
   FA_X1 i_61 (.A(n_116), .B(n_114), .CI(n_112), .CO(n_123), .S(n_122));
   FA_X1 i_62 (.A(n_110), .B(n_120), .CI(n_118), .CO(n_125), .S(n_124));
   FA_X1 i_63 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_64 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   HA_X1 i_65 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_66 (.A(n_485), .B(n_487), .CI(n_498), .CO(n_133), .S(n_132));
   FA_X1 i_67 (.A(n_511), .B(n_524), .CI(n_535), .CO(n_135), .S(n_134));
   FA_X1 i_68 (.A(n_547), .B(n_560), .CI(n_571), .CO(n_137), .S(n_136));
   FA_X1 i_69 (.A(n_583), .B(n_595), .CI(n_606), .CO(n_139), .S(n_138));
   FA_X1 i_70 (.A(n_619), .B(n_630), .CI(n_117), .CO(n_141), .S(n_140));
   FA_X1 i_71 (.A(n_115), .B(n_113), .CI(n_111), .CO(n_143), .S(n_142));
   FA_X1 i_72 (.A(n_119), .B(n_140), .CI(n_138), .CO(n_145), .S(n_144));
   FA_X1 i_73 (.A(n_136), .B(n_134), .CI(n_132), .CO(n_147), .S(n_146));
   FA_X1 i_74 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_75 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_76 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_77 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   FA_X1 i_78 (.A(n_497), .B(n_510), .CI(n_523), .CO(n_157), .S(n_156));
   FA_X1 i_79 (.A(n_534), .B(n_546), .CI(n_559), .CO(n_159), .S(n_158));
   FA_X1 i_80 (.A(n_570), .B(n_582), .CI(n_594), .CO(n_161), .S(n_160));
   FA_X1 i_81 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_163), .S(n_162));
   FA_X1 i_82 (.A(n_133), .B(n_143), .CI(n_141), .CO(n_165), .S(n_164));
   FA_X1 i_83 (.A(n_471), .B(n_160), .CI(n_158), .CO(n_167), .S(n_166));
   FA_X1 i_84 (.A(n_156), .B(n_479), .CI(n_162), .CO(n_169), .S(n_168));
   FA_X1 i_85 (.A(n_147), .B(n_145), .CI(n_164), .CO(n_171), .S(n_170));
   FA_X1 i_86 (.A(n_149), .B(n_168), .CI(n_166), .CO(n_173), .S(n_172));
   FA_X1 i_87 (.A(n_170), .B(n_151), .CI(n_172), .CO(n_175), .S(n_174));
   HA_X1 i_88 (.A(n_153), .B(n_155), .CO(n_177), .S(n_176));
   FA_X1 i_89 (.A(n_486), .B(n_496), .CI(n_509), .CO(n_179), .S(n_178));
   FA_X1 i_90 (.A(n_522), .B(n_533), .CI(n_545), .CO(n_181), .S(n_180));
   FA_X1 i_91 (.A(n_558), .B(n_569), .CI(n_581), .CO(n_183), .S(n_182));
   FA_X1 i_92 (.A(n_470), .B(n_161), .CI(n_159), .CO(n_185), .S(n_184));
   FA_X1 i_93 (.A(n_157), .B(n_477), .CI(n_163), .CO(n_187), .S(n_186));
   FA_X1 i_94 (.A(n_460), .B(n_182), .CI(n_180), .CO(n_189), .S(n_188));
   FA_X1 i_95 (.A(n_178), .B(n_466), .CI(n_165), .CO(n_191), .S(n_190));
   FA_X1 i_96 (.A(n_186), .B(n_184), .CI(n_167), .CO(n_193), .S(n_192));
   FA_X1 i_97 (.A(n_169), .B(n_190), .CI(n_188), .CO(n_195), .S(n_194));
   FA_X1 i_98 (.A(n_171), .B(n_192), .CI(n_173), .CO(n_197), .S(n_196));
   FA_X1 i_99 (.A(n_194), .B(n_196), .CI(n_175), .CO(n_199), .S(n_198));
   FA_X1 i_100 (.A(n_495), .B(n_508), .CI(n_521), .CO(n_201), .S(n_200));
   FA_X1 i_101 (.A(n_532), .B(n_544), .CI(n_557), .CO(n_203), .S(n_202));
   FA_X1 i_102 (.A(n_568), .B(n_580), .CI(n_593), .CO(n_205), .S(n_204));
   FA_X1 i_103 (.A(n_181), .B(n_179), .CI(n_467), .CO(n_207), .S(n_206));
   FA_X1 i_104 (.A(n_185), .B(n_204), .CI(n_202), .CO(n_209), .S(n_208));
   FA_X1 i_105 (.A(n_200), .B(n_454), .CI(n_187), .CO(n_211), .S(n_210));
   FA_X1 i_106 (.A(n_206), .B(n_445), .CI(n_189), .CO(n_213), .S(n_212));
   FA_X1 i_107 (.A(n_191), .B(n_193), .CI(n_210), .CO(n_215), .S(n_214));
   FA_X1 i_108 (.A(n_208), .B(n_212), .CI(n_195), .CO(n_217), .S(n_216));
   FA_X1 i_109 (.A(n_214), .B(n_197), .CI(n_216), .CO(n_219), .S(n_218));
   FA_X1 i_110 (.A(n_494), .B(n_507), .CI(n_520), .CO(n_221), .S(n_220));
   FA_X1 i_111 (.A(n_531), .B(n_543), .CI(n_556), .CO(n_223), .S(n_222));
   FA_X1 i_112 (.A(n_205), .B(n_203), .CI(n_201), .CO(n_225), .S(n_224));
   FA_X1 i_113 (.A(n_452), .B(n_207), .CI(n_447), .CO(n_227), .S(n_226));
   FA_X1 i_114 (.A(n_430), .B(n_222), .CI(n_220), .CO(n_229), .S(n_228));
   FA_X1 i_115 (.A(n_439), .B(n_224), .CI(n_209), .CO(n_231), .S(n_230));
   FA_X1 i_116 (.A(n_211), .B(n_226), .CI(n_213), .CO(n_233), .S(n_232));
   FA_X1 i_117 (.A(n_228), .B(n_230), .CI(n_215), .CO(n_235), .S(n_234));
   FA_X1 i_118 (.A(n_232), .B(n_217), .CI(n_234), .CO(n_237), .S(n_236));
   FA_X1 i_119 (.A(n_493), .B(n_506), .CI(n_519), .CO(n_239), .S(n_238));
   FA_X1 i_120 (.A(n_530), .B(n_542), .CI(n_555), .CO(n_241), .S(n_240));
   FA_X1 i_121 (.A(n_223), .B(n_221), .CI(n_437), .CO(n_243), .S(n_242));
   FA_X1 i_122 (.A(n_225), .B(n_416), .CI(n_240), .CO(n_245), .S(n_244));
   FA_X1 i_123 (.A(n_238), .B(n_424), .CI(n_227), .CO(n_247), .S(n_246));
   FA_X1 i_124 (.A(n_242), .B(n_229), .CI(n_231), .CO(n_249), .S(n_248));
   FA_X1 i_125 (.A(n_246), .B(n_244), .CI(n_233), .CO(n_251), .S(n_250));
   FA_X1 i_126 (.A(n_248), .B(n_235), .CI(n_250), .CO(n_253), .S(n_252));
   FA_X1 i_127 (.A(n_492), .B(n_505), .CI(n_518), .CO(n_255), .S(n_254));
   FA_X1 i_128 (.A(n_529), .B(n_541), .CI(n_554), .CO(n_257), .S(n_256));
   FA_X1 i_129 (.A(n_422), .B(n_243), .CI(n_415), .CO(n_259), .S(n_258));
   FA_X1 i_130 (.A(n_256), .B(n_254), .CI(n_409), .CO(n_261), .S(n_260));
   FA_X1 i_131 (.A(n_402), .B(n_245), .CI(n_247), .CO(n_263), .S(n_262));
   FA_X1 i_132 (.A(n_258), .B(n_260), .CI(n_249), .CO(n_265), .S(n_264));
   FA_X1 i_133 (.A(n_262), .B(n_251), .CI(n_264), .CO(n_267), .S(n_266));
   FA_X1 i_134 (.A(n_491), .B(n_504), .CI(n_517), .CO(n_269), .S(n_268));
   FA_X1 i_135 (.A(n_257), .B(n_255), .CI(n_407), .CO(n_271), .S(n_270));
   FA_X1 i_136 (.A(n_400), .B(n_385), .CI(n_268), .CO(n_273), .S(n_272));
   FA_X1 i_137 (.A(n_394), .B(n_259), .CI(n_270), .CO(n_275), .S(n_274));
   FA_X1 i_138 (.A(n_261), .B(n_263), .CI(n_272), .CO(n_277), .S(n_276));
   FA_X1 i_139 (.A(n_274), .B(n_265), .CI(n_276), .CO(n_279), .S(n_278));
   FA_X1 i_140 (.A(n_490), .B(n_503), .CI(n_516), .CO(n_281), .S(n_280));
   FA_X1 i_141 (.A(n_269), .B(n_392), .CI(n_271), .CO(n_283), .S(n_282));
   FA_X1 i_142 (.A(n_372), .B(n_280), .CI(n_378), .CO(n_285), .S(n_284));
   FA_X1 i_143 (.A(n_282), .B(n_273), .CI(n_275), .CO(n_287), .S(n_286));
   FA_X1 i_144 (.A(n_284), .B(n_286), .CI(n_277), .CO(n_289), .S(n_288));
   FA_X1 i_145 (.A(n_489), .B(n_502), .CI(n_515), .CO(n_291), .S(n_290));
   FA_X1 i_146 (.A(n_371), .B(n_290), .CI(n_365), .CO(n_293), .S(n_292));
   FA_X1 i_147 (.A(n_283), .B(n_357), .CI(n_285), .CO(n_295), .S(n_294));
   FA_X1 i_148 (.A(n_292), .B(n_287), .CI(n_294), .CO(n_297), .S(n_296));
   FA_X1 i_149 (.A(n_291), .B(n_363), .CI(n_356), .CO(n_299), .S(n_298));
   FA_X1 i_150 (.A(n_342), .B(n_350), .CI(n_298), .CO(n_301), .S(n_300));
   FA_X1 i_151 (.A(n_293), .B(n_295), .CI(n_300), .CO(n_303), .S(n_302));
   FA_X1 i_152 (.A(n_348), .B(n_329), .CI(n_335), .CO(n_305), .S(n_304));
   FA_X1 i_153 (.A(n_299), .B(n_301), .CI(n_304), .CO(n_307), .S(n_306));
   FA_X1 i_154 (.A(n_323), .B(n_315), .CI(n_305), .CO(n_309), .S(n_308));
   FA_X1 i_155 (.A(n_321), .B(n_312), .CI(n_314), .CO(n_311), .S(n_310));
   XOR2_X1 i_156 (.A(n_796), .B(n_313), .Z(n_312));
   NOR2_X1 i_157 (.A1(n_799), .A2(n_798), .ZN(n_313));
   OAI22_X1 i_158 (.A1(n_320), .A2(n_319), .B1(n_318), .B2(n_316), .ZN(n_314));
   XNOR2_X1 i_159 (.A(n_317), .B(n_316), .ZN(n_315));
   OAI22_X1 i_160 (.A1(n_340), .A2(n_339), .B1(n_341), .B2(n_337), .ZN(n_316));
   XOR2_X1 i_161 (.A(n_320), .B(n_319), .Z(n_317));
   AND2_X1 i_162 (.A1(n_320), .A2(n_319), .ZN(n_318));
   OAI22_X1 i_163 (.A1(n_347), .A2(n_333), .B1(n_332), .B2(n_330), .ZN(n_319));
   NOR2_X1 i_164 (.A1(n_834), .A2(n_822), .ZN(n_320));
   NAND2_X1 i_165 (.A1(n_325), .A2(n_322), .ZN(n_321));
   OAI21_X1 i_166 (.A(n_328), .B1(n_327), .B2(n_326), .ZN(n_322));
   XNOR2_X1 i_167 (.A(n_328), .B(n_324), .ZN(n_323));
   OAI21_X1 i_168 (.A(n_325), .B1(n_327), .B2(n_326), .ZN(n_324));
   NAND2_X1 i_169 (.A1(n_327), .A2(n_326), .ZN(n_325));
   NOR2_X1 i_170 (.A1(n_836), .A2(n_820), .ZN(n_326));
   NAND2_X1 i_171 (.A1(operand2[14]), .A2(operand1[11]), .ZN(n_327));
   NOR2_X1 i_172 (.A1(n_835), .A2(n_821), .ZN(n_328));
   XOR2_X1 i_173 (.A(n_331), .B(n_330), .Z(n_329));
   OAI22_X1 i_174 (.A1(n_501), .A2(n_346), .B1(n_345), .B2(n_343), .ZN(n_330));
   AOI21_X1 i_175 (.A(n_332), .B1(n_346), .B2(n_334), .ZN(n_331));
   NOR2_X1 i_176 (.A1(n_346), .A2(n_334), .ZN(n_332));
   INV_X1 i_177 (.A(n_334), .ZN(n_333));
   NOR2_X1 i_178 (.A1(n_833), .A2(n_822), .ZN(n_334));
   XNOR2_X1 i_179 (.A(n_341), .B(n_336), .ZN(n_335));
   OAI21_X1 i_180 (.A(n_338), .B1(n_340), .B2(n_339), .ZN(n_336));
   INV_X1 i_181 (.A(n_338), .ZN(n_337));
   NAND2_X1 i_182 (.A1(n_340), .A2(n_339), .ZN(n_338));
   NOR2_X1 i_183 (.A1(n_836), .A2(n_819), .ZN(n_339));
   NAND2_X1 i_184 (.A1(operand2[14]), .A2(operand1[10]), .ZN(n_340));
   NOR2_X1 i_185 (.A1(n_835), .A2(n_820), .ZN(n_341));
   XNOR2_X1 i_186 (.A(n_344), .B(n_343), .ZN(n_342));
   NOR2_X1 i_187 (.A1(n_832), .A2(n_822), .ZN(n_343));
   AOI21_X1 i_188 (.A(n_345), .B1(n_502), .B2(n_347), .ZN(n_344));
   AOI22_X1 i_189 (.A1(operand2[11]), .A2(operand1[12]), .B1(operand2[10]), 
      .B2(operand1[13]), .ZN(n_345));
   INV_X1 i_190 (.A(n_347), .ZN(n_346));
   NOR2_X1 i_191 (.A1(n_834), .A2(n_821), .ZN(n_347));
   NAND2_X1 i_192 (.A1(n_352), .A2(n_349), .ZN(n_348));
   OAI21_X1 i_193 (.A(n_355), .B1(n_354), .B2(n_353), .ZN(n_349));
   XNOR2_X1 i_194 (.A(n_355), .B(n_351), .ZN(n_350));
   OAI21_X1 i_195 (.A(n_352), .B1(n_354), .B2(n_353), .ZN(n_351));
   NAND2_X1 i_196 (.A1(n_354), .A2(n_353), .ZN(n_352));
   NOR2_X1 i_197 (.A1(n_836), .A2(n_818), .ZN(n_353));
   NAND2_X1 i_198 (.A1(operand2[14]), .A2(operand1[9]), .ZN(n_354));
   NOR2_X1 i_199 (.A1(n_835), .A2(n_819), .ZN(n_355));
   OAI21_X1 i_200 (.A(n_361), .B1(n_360), .B2(n_358), .ZN(n_356));
   XNOR2_X1 i_201 (.A(n_359), .B(n_358), .ZN(n_357));
   OAI22_X1 i_202 (.A1(n_383), .A2(n_382), .B1(n_384), .B2(n_380), .ZN(n_358));
   AOI21_X1 i_203 (.A(n_360), .B1(n_281), .B2(n_362), .ZN(n_359));
   NOR2_X1 i_204 (.A1(n_281), .A2(n_362), .ZN(n_360));
   NAND2_X1 i_205 (.A1(n_281), .A2(n_362), .ZN(n_361));
   NAND2_X1 i_206 (.A1(operand2[8]), .A2(operand1[14]), .ZN(n_362));
   NAND2_X1 i_207 (.A1(n_367), .A2(n_364), .ZN(n_363));
   OAI21_X1 i_208 (.A(n_370), .B1(n_369), .B2(n_368), .ZN(n_364));
   XNOR2_X1 i_209 (.A(n_370), .B(n_366), .ZN(n_365));
   OAI21_X1 i_210 (.A(n_367), .B1(n_369), .B2(n_368), .ZN(n_366));
   NAND2_X1 i_211 (.A1(n_369), .A2(n_368), .ZN(n_367));
   NOR2_X1 i_212 (.A1(n_836), .A2(n_817), .ZN(n_368));
   NAND2_X1 i_213 (.A1(operand2[14]), .A2(operand1[8]), .ZN(n_369));
   NOR2_X1 i_214 (.A1(n_835), .A2(n_818), .ZN(n_370));
   OAI22_X1 i_215 (.A1(n_391), .A2(n_377), .B1(n_375), .B2(n_373), .ZN(n_371));
   XOR2_X1 i_216 (.A(n_374), .B(n_373), .Z(n_372));
   NOR2_X1 i_217 (.A1(n_390), .A2(n_386), .ZN(n_373));
   OAI21_X1 i_218 (.A(n_376), .B1(n_391), .B2(n_377), .ZN(n_374));
   INV_X1 i_219 (.A(n_376), .ZN(n_375));
   NAND2_X1 i_220 (.A1(n_391), .A2(n_377), .ZN(n_376));
   NOR2_X1 i_221 (.A1(n_830), .A2(n_822), .ZN(n_377));
   XNOR2_X1 i_222 (.A(n_384), .B(n_379), .ZN(n_378));
   OAI21_X1 i_223 (.A(n_381), .B1(n_383), .B2(n_382), .ZN(n_379));
   INV_X1 i_224 (.A(n_381), .ZN(n_380));
   NAND2_X1 i_225 (.A1(n_383), .A2(n_382), .ZN(n_381));
   NOR2_X1 i_226 (.A1(n_836), .A2(n_816), .ZN(n_382));
   NAND2_X1 i_227 (.A1(operand2[14]), .A2(operand1[7]), .ZN(n_383));
   NOR2_X1 i_228 (.A1(n_835), .A2(n_817), .ZN(n_384));
   XNOR2_X1 i_229 (.A(n_388), .B(n_387), .ZN(n_385));
   NOR2_X1 i_230 (.A1(n_389), .A2(n_387), .ZN(n_386));
   NOR2_X1 i_231 (.A1(n_829), .A2(n_822), .ZN(n_387));
   NOR2_X1 i_232 (.A1(n_390), .A2(n_389), .ZN(n_388));
   AOI22_X1 i_233 (.A1(operand2[8]), .A2(operand1[12]), .B1(operand2[7]), 
      .B2(operand1[13]), .ZN(n_389));
   NOR3_X1 i_234 (.A1(n_830), .A2(n_820), .A3(n_391), .ZN(n_390));
   NAND2_X1 i_235 (.A1(operand2[8]), .A2(operand1[13]), .ZN(n_391));
   NAND2_X1 i_236 (.A1(n_396), .A2(n_393), .ZN(n_392));
   OAI21_X1 i_237 (.A(n_399), .B1(n_398), .B2(n_397), .ZN(n_393));
   XNOR2_X1 i_238 (.A(n_399), .B(n_395), .ZN(n_394));
   OAI21_X1 i_239 (.A(n_396), .B1(n_398), .B2(n_397), .ZN(n_395));
   NAND2_X1 i_240 (.A1(n_398), .A2(n_397), .ZN(n_396));
   NOR2_X1 i_241 (.A1(n_836), .A2(n_815), .ZN(n_397));
   NAND2_X1 i_242 (.A1(operand2[14]), .A2(operand1[6]), .ZN(n_398));
   NOR2_X1 i_243 (.A1(n_835), .A2(n_816), .ZN(n_399));
   NOR2_X1 i_244 (.A1(n_404), .A2(n_401), .ZN(n_400));
   NOR2_X1 i_245 (.A1(n_241), .A2(n_405), .ZN(n_401));
   XOR2_X1 i_246 (.A(n_241), .B(n_403), .Z(n_402));
   NOR2_X1 i_247 (.A1(n_405), .A2(n_404), .ZN(n_403));
   NOR2_X1 i_248 (.A1(n_239), .A2(n_406), .ZN(n_404));
   AND2_X1 i_249 (.A1(n_239), .A2(n_406), .ZN(n_405));
   NAND2_X1 i_250 (.A1(operand2[5]), .A2(operand1[14]), .ZN(n_406));
   NAND2_X1 i_251 (.A1(n_411), .A2(n_408), .ZN(n_407));
   OAI21_X1 i_252 (.A(n_414), .B1(n_413), .B2(n_412), .ZN(n_408));
   XNOR2_X1 i_253 (.A(n_414), .B(n_410), .ZN(n_409));
   OAI21_X1 i_254 (.A(n_411), .B1(n_413), .B2(n_412), .ZN(n_410));
   NAND2_X1 i_255 (.A1(n_413), .A2(n_412), .ZN(n_411));
   NOR2_X1 i_256 (.A1(n_836), .A2(n_814), .ZN(n_412));
   NAND2_X1 i_257 (.A1(operand2[14]), .A2(operand1[5]), .ZN(n_413));
   NOR2_X1 i_258 (.A1(n_835), .A2(n_815), .ZN(n_414));
   OAI22_X1 i_259 (.A1(n_436), .A2(n_421), .B1(n_419), .B2(n_417), .ZN(n_415));
   XOR2_X1 i_260 (.A(n_418), .B(n_417), .Z(n_416));
   NOR2_X1 i_261 (.A1(n_435), .A2(n_431), .ZN(n_417));
   OAI21_X1 i_262 (.A(n_420), .B1(n_436), .B2(n_421), .ZN(n_418));
   INV_X1 i_263 (.A(n_420), .ZN(n_419));
   NAND2_X1 i_264 (.A1(n_436), .A2(n_421), .ZN(n_420));
   NOR2_X1 i_265 (.A1(n_827), .A2(n_822), .ZN(n_421));
   NAND2_X1 i_266 (.A1(n_426), .A2(n_423), .ZN(n_422));
   OAI21_X1 i_267 (.A(n_429), .B1(n_428), .B2(n_427), .ZN(n_423));
   XNOR2_X1 i_268 (.A(n_429), .B(n_425), .ZN(n_424));
   OAI21_X1 i_269 (.A(n_426), .B1(n_428), .B2(n_427), .ZN(n_425));
   NAND2_X1 i_270 (.A1(n_428), .A2(n_427), .ZN(n_426));
   NOR2_X1 i_271 (.A1(n_836), .A2(n_813), .ZN(n_427));
   NAND2_X1 i_272 (.A1(operand2[14]), .A2(operand1[4]), .ZN(n_428));
   NOR2_X1 i_273 (.A1(n_835), .A2(n_814), .ZN(n_429));
   XNOR2_X1 i_274 (.A(n_433), .B(n_432), .ZN(n_430));
   NOR2_X1 i_275 (.A1(n_434), .A2(n_432), .ZN(n_431));
   NOR2_X1 i_276 (.A1(n_826), .A2(n_822), .ZN(n_432));
   NOR2_X1 i_277 (.A1(n_435), .A2(n_434), .ZN(n_433));
   AOI22_X1 i_278 (.A1(operand2[5]), .A2(operand1[12]), .B1(operand2[4]), 
      .B2(operand1[13]), .ZN(n_434));
   NOR3_X1 i_279 (.A1(n_827), .A2(n_820), .A3(n_436), .ZN(n_435));
   NAND2_X1 i_280 (.A1(operand2[5]), .A2(operand1[13]), .ZN(n_436));
   NAND2_X1 i_281 (.A1(n_441), .A2(n_438), .ZN(n_437));
   OAI21_X1 i_282 (.A(n_444), .B1(n_443), .B2(n_442), .ZN(n_438));
   XNOR2_X1 i_283 (.A(n_444), .B(n_440), .ZN(n_439));
   OAI21_X1 i_284 (.A(n_441), .B1(n_443), .B2(n_442), .ZN(n_440));
   NAND2_X1 i_285 (.A1(n_443), .A2(n_442), .ZN(n_441));
   NOR2_X1 i_286 (.A1(n_836), .A2(n_812), .ZN(n_442));
   NAND2_X1 i_287 (.A1(operand2[14]), .A2(operand1[3]), .ZN(n_443));
   NOR2_X1 i_288 (.A1(n_835), .A2(n_813), .ZN(n_444));
   AOI22_X1 i_289 (.A1(n_449), .A2(n_447), .B1(n_807), .B2(n_446), .ZN(n_445));
   OAI21_X1 i_290 (.A(n_449), .B1(n_451), .B2(n_450), .ZN(n_446));
   OAI21_X1 i_291 (.A(n_449), .B1(n_807), .B2(n_448), .ZN(n_447));
   NOR2_X1 i_292 (.A1(n_451), .A2(n_450), .ZN(n_448));
   NAND2_X1 i_293 (.A1(n_451), .A2(n_450), .ZN(n_449));
   OAI21_X1 i_294 (.A(n_464), .B1(n_463), .B2(n_461), .ZN(n_450));
   NAND2_X1 i_295 (.A1(operand2[2]), .A2(operand1[14]), .ZN(n_451));
   NAND2_X1 i_296 (.A1(n_456), .A2(n_453), .ZN(n_452));
   OAI21_X1 i_297 (.A(n_459), .B1(n_458), .B2(n_457), .ZN(n_453));
   XNOR2_X1 i_298 (.A(n_459), .B(n_455), .ZN(n_454));
   OAI21_X1 i_299 (.A(n_456), .B1(n_458), .B2(n_457), .ZN(n_455));
   NAND2_X1 i_300 (.A1(n_458), .A2(n_457), .ZN(n_456));
   NOR2_X1 i_301 (.A1(n_836), .A2(n_811), .ZN(n_457));
   NAND2_X1 i_302 (.A1(operand2[14]), .A2(operand1[2]), .ZN(n_458));
   NOR2_X1 i_303 (.A1(n_835), .A2(n_812), .ZN(n_459));
   XNOR2_X1 i_304 (.A(n_462), .B(n_461), .ZN(n_460));
   NOR2_X1 i_305 (.A1(n_824), .A2(n_822), .ZN(n_461));
   NOR2_X1 i_306 (.A1(n_465), .A2(n_463), .ZN(n_462));
   AOI21_X1 i_307 (.A(n_476), .B1(operand2[3]), .B2(operand1[12]), .ZN(n_463));
   INV_X1 i_308 (.A(n_465), .ZN(n_464));
   NOR3_X1 i_309 (.A1(n_826), .A2(n_820), .A3(n_475), .ZN(n_465));
   OAI21_X1 i_310 (.A(n_467), .B1(n_469), .B2(n_468), .ZN(n_466));
   NAND2_X1 i_311 (.A1(n_469), .A2(n_468), .ZN(n_467));
   NAND2_X1 i_312 (.A1(operand2[13]), .A2(operand1[2]), .ZN(n_468));
   NOR2_X1 i_313 (.A1(n_837), .A2(n_809), .ZN(n_469));
   OAI22_X1 i_314 (.A1(n_618), .A2(n_475), .B1(n_474), .B2(n_472), .ZN(n_470));
   XNOR2_X1 i_315 (.A(n_473), .B(n_472), .ZN(n_471));
   NOR2_X1 i_316 (.A1(n_823), .A2(n_822), .ZN(n_472));
   AOI21_X1 i_317 (.A(n_474), .B1(n_619), .B2(n_476), .ZN(n_473));
   AOI22_X1 i_318 (.A1(operand2[2]), .A2(operand1[12]), .B1(operand2[1]), 
      .B2(operand1[13]), .ZN(n_474));
   INV_X1 i_319 (.A(n_476), .ZN(n_475));
   NOR2_X1 i_320 (.A1(n_825), .A2(n_821), .ZN(n_476));
   NAND2_X1 i_321 (.A1(n_481), .A2(n_478), .ZN(n_477));
   OAI21_X1 i_322 (.A(n_484), .B1(n_483), .B2(n_482), .ZN(n_478));
   XNOR2_X1 i_323 (.A(n_484), .B(n_480), .ZN(n_479));
   OAI21_X1 i_324 (.A(n_481), .B1(n_483), .B2(n_482), .ZN(n_480));
   NAND2_X1 i_325 (.A1(n_483), .A2(n_482), .ZN(n_481));
   NOR2_X1 i_326 (.A1(n_836), .A2(n_809), .ZN(n_482));
   NAND2_X1 i_327 (.A1(operand2[14]), .A2(operand1[0]), .ZN(n_483));
   NOR2_X1 i_328 (.A1(n_835), .A2(n_810), .ZN(n_484));
   NOR2_X1 i_329 (.A1(n_836), .A2(n_808), .ZN(n_485));
   NOR2_X1 i_330 (.A1(n_835), .A2(n_811), .ZN(n_486));
   NOR2_X1 i_331 (.A1(n_835), .A2(n_809), .ZN(n_487));
   NOR2_X1 i_332 (.A1(n_835), .A2(n_808), .ZN(n_488));
   NOR2_X1 i_333 (.A1(n_834), .A2(n_819), .ZN(n_489));
   NOR2_X1 i_334 (.A1(n_834), .A2(n_818), .ZN(n_490));
   NOR2_X1 i_335 (.A1(n_834), .A2(n_817), .ZN(n_491));
   NOR2_X1 i_336 (.A1(n_834), .A2(n_816), .ZN(n_492));
   NOR2_X1 i_337 (.A1(n_834), .A2(n_815), .ZN(n_493));
   NOR2_X1 i_338 (.A1(n_834), .A2(n_814), .ZN(n_494));
   NOR2_X1 i_339 (.A1(n_834), .A2(n_813), .ZN(n_495));
   NOR2_X1 i_340 (.A1(n_834), .A2(n_812), .ZN(n_496));
   NOR2_X1 i_341 (.A1(n_834), .A2(n_811), .ZN(n_497));
   NOR2_X1 i_342 (.A1(n_834), .A2(n_810), .ZN(n_498));
   NOR2_X1 i_343 (.A1(n_834), .A2(n_809), .ZN(n_499));
   NOR2_X1 i_344 (.A1(n_834), .A2(n_808), .ZN(n_500));
   INV_X1 i_345 (.A(n_502), .ZN(n_501));
   NOR2_X1 i_346 (.A1(n_833), .A2(n_820), .ZN(n_502));
   NOR2_X1 i_347 (.A1(n_833), .A2(n_819), .ZN(n_503));
   NOR2_X1 i_348 (.A1(n_833), .A2(n_818), .ZN(n_504));
   NOR2_X1 i_349 (.A1(n_833), .A2(n_817), .ZN(n_505));
   NOR2_X1 i_350 (.A1(n_833), .A2(n_816), .ZN(n_506));
   NOR2_X1 i_351 (.A1(n_833), .A2(n_815), .ZN(n_507));
   NOR2_X1 i_352 (.A1(n_833), .A2(n_814), .ZN(n_508));
   NOR2_X1 i_353 (.A1(n_833), .A2(n_813), .ZN(n_509));
   NOR2_X1 i_354 (.A1(n_833), .A2(n_812), .ZN(n_510));
   NOR2_X1 i_355 (.A1(n_833), .A2(n_811), .ZN(n_511));
   NOR2_X1 i_356 (.A1(n_833), .A2(n_810), .ZN(n_512));
   NOR2_X1 i_357 (.A1(n_833), .A2(n_809), .ZN(n_513));
   NOR2_X1 i_358 (.A1(n_833), .A2(n_808), .ZN(n_514));
   NOR2_X1 i_359 (.A1(n_832), .A2(n_821), .ZN(n_515));
   NOR2_X1 i_360 (.A1(n_832), .A2(n_820), .ZN(n_516));
   NOR2_X1 i_361 (.A1(n_832), .A2(n_819), .ZN(n_517));
   NOR2_X1 i_362 (.A1(n_832), .A2(n_818), .ZN(n_518));
   NOR2_X1 i_363 (.A1(n_832), .A2(n_817), .ZN(n_519));
   NOR2_X1 i_364 (.A1(n_832), .A2(n_816), .ZN(n_520));
   NOR2_X1 i_365 (.A1(n_832), .A2(n_815), .ZN(n_521));
   NOR2_X1 i_366 (.A1(n_832), .A2(n_814), .ZN(n_522));
   NOR2_X1 i_367 (.A1(n_832), .A2(n_813), .ZN(n_523));
   NOR2_X1 i_368 (.A1(n_832), .A2(n_812), .ZN(n_524));
   NOR2_X1 i_369 (.A1(n_832), .A2(n_811), .ZN(n_525));
   NOR2_X1 i_370 (.A1(n_832), .A2(n_810), .ZN(n_526));
   NOR2_X1 i_371 (.A1(n_832), .A2(n_809), .ZN(n_527));
   NOR2_X1 i_372 (.A1(n_832), .A2(n_808), .ZN(n_528));
   NOR2_X1 i_373 (.A1(n_831), .A2(n_819), .ZN(n_529));
   NOR2_X1 i_374 (.A1(n_831), .A2(n_818), .ZN(n_530));
   NOR2_X1 i_375 (.A1(n_831), .A2(n_817), .ZN(n_531));
   NOR2_X1 i_376 (.A1(n_831), .A2(n_816), .ZN(n_532));
   NOR2_X1 i_377 (.A1(n_831), .A2(n_815), .ZN(n_533));
   NOR2_X1 i_378 (.A1(n_831), .A2(n_814), .ZN(n_534));
   NOR2_X1 i_379 (.A1(n_831), .A2(n_813), .ZN(n_535));
   NOR2_X1 i_380 (.A1(n_831), .A2(n_812), .ZN(n_536));
   NOR2_X1 i_381 (.A1(n_831), .A2(n_811), .ZN(n_537));
   NOR2_X1 i_382 (.A1(n_831), .A2(n_810), .ZN(n_538));
   NOR2_X1 i_383 (.A1(n_831), .A2(n_809), .ZN(n_539));
   NOR2_X1 i_384 (.A1(n_831), .A2(n_808), .ZN(n_540));
   NOR2_X1 i_385 (.A1(n_830), .A2(n_820), .ZN(n_541));
   NOR2_X1 i_386 (.A1(n_830), .A2(n_819), .ZN(n_542));
   NOR2_X1 i_387 (.A1(n_830), .A2(n_818), .ZN(n_543));
   NOR2_X1 i_388 (.A1(n_830), .A2(n_817), .ZN(n_544));
   NOR2_X1 i_389 (.A1(n_830), .A2(n_816), .ZN(n_545));
   NOR2_X1 i_390 (.A1(n_830), .A2(n_815), .ZN(n_546));
   NOR2_X1 i_391 (.A1(n_830), .A2(n_814), .ZN(n_547));
   NOR2_X1 i_392 (.A1(n_830), .A2(n_813), .ZN(n_548));
   NOR2_X1 i_393 (.A1(n_830), .A2(n_812), .ZN(n_549));
   NOR2_X1 i_394 (.A1(n_830), .A2(n_811), .ZN(n_550));
   NOR2_X1 i_395 (.A1(n_830), .A2(n_810), .ZN(n_551));
   NOR2_X1 i_396 (.A1(n_830), .A2(n_809), .ZN(n_552));
   NOR2_X1 i_397 (.A1(n_830), .A2(n_808), .ZN(n_553));
   NOR2_X1 i_398 (.A1(n_829), .A2(n_821), .ZN(n_554));
   NOR2_X1 i_399 (.A1(n_829), .A2(n_820), .ZN(n_555));
   NOR2_X1 i_400 (.A1(n_829), .A2(n_819), .ZN(n_556));
   NOR2_X1 i_401 (.A1(n_829), .A2(n_818), .ZN(n_557));
   NOR2_X1 i_402 (.A1(n_829), .A2(n_817), .ZN(n_558));
   NOR2_X1 i_403 (.A1(n_829), .A2(n_816), .ZN(n_559));
   NOR2_X1 i_404 (.A1(n_829), .A2(n_815), .ZN(n_560));
   NOR2_X1 i_405 (.A1(n_829), .A2(n_814), .ZN(n_561));
   NOR2_X1 i_406 (.A1(n_829), .A2(n_813), .ZN(n_562));
   NOR2_X1 i_407 (.A1(n_829), .A2(n_812), .ZN(n_563));
   NOR2_X1 i_408 (.A1(n_829), .A2(n_811), .ZN(n_564));
   NOR2_X1 i_409 (.A1(n_829), .A2(n_810), .ZN(n_565));
   NOR2_X1 i_410 (.A1(n_829), .A2(n_809), .ZN(n_566));
   NOR2_X1 i_411 (.A1(n_829), .A2(n_808), .ZN(n_567));
   NOR2_X1 i_412 (.A1(n_828), .A2(n_819), .ZN(n_568));
   NOR2_X1 i_413 (.A1(n_828), .A2(n_818), .ZN(n_569));
   NOR2_X1 i_414 (.A1(n_828), .A2(n_817), .ZN(n_570));
   NOR2_X1 i_415 (.A1(n_828), .A2(n_816), .ZN(n_571));
   NOR2_X1 i_416 (.A1(n_828), .A2(n_815), .ZN(n_572));
   NOR2_X1 i_417 (.A1(n_828), .A2(n_814), .ZN(n_573));
   NOR2_X1 i_418 (.A1(n_828), .A2(n_813), .ZN(n_574));
   NOR2_X1 i_419 (.A1(n_828), .A2(n_812), .ZN(n_575));
   NOR2_X1 i_421 (.A1(n_828), .A2(n_810), .ZN(n_577));
   NOR2_X1 i_422 (.A1(n_828), .A2(n_809), .ZN(n_578));
   NOR2_X1 i_424 (.A1(n_827), .A2(n_820), .ZN(n_580));
   NOR2_X1 i_425 (.A1(n_827), .A2(n_819), .ZN(n_581));
   NOR2_X1 i_426 (.A1(n_827), .A2(n_818), .ZN(n_582));
   NOR2_X1 i_427 (.A1(n_827), .A2(n_817), .ZN(n_583));
   NOR2_X1 i_428 (.A1(n_827), .A2(n_816), .ZN(n_584));
   NOR2_X1 i_429 (.A1(n_827), .A2(n_815), .ZN(n_585));
   NOR2_X1 i_430 (.A1(n_827), .A2(n_814), .ZN(n_586));
   NOR2_X1 i_431 (.A1(n_827), .A2(n_813), .ZN(n_587));
   NOR2_X1 i_433 (.A1(n_827), .A2(n_811), .ZN(n_589));
   NOR2_X1 i_434 (.A1(n_827), .A2(n_810), .ZN(n_590));
   NOR2_X1 i_436 (.A1(n_827), .A2(n_808), .ZN(n_592));
   NOR2_X1 i_437 (.A1(n_826), .A2(n_821), .ZN(n_593));
   NOR2_X1 i_438 (.A1(n_826), .A2(n_819), .ZN(n_594));
   NOR2_X1 i_439 (.A1(n_826), .A2(n_818), .ZN(n_595));
   NOR2_X1 i_440 (.A1(n_826), .A2(n_817), .ZN(n_596));
   NOR2_X1 i_441 (.A1(n_826), .A2(n_816), .ZN(n_597));
   NOR2_X1 i_442 (.A1(n_826), .A2(n_815), .ZN(n_598));
   NOR2_X1 i_443 (.A1(n_826), .A2(n_814), .ZN(n_599));
   NOR2_X1 i_445 (.A1(n_826), .A2(n_812), .ZN(n_601));
   NOR2_X1 i_448 (.A1(n_826), .A2(n_809), .ZN(n_604));
   NOR2_X1 i_449 (.A1(n_826), .A2(n_808), .ZN(n_605));
   NOR2_X1 i_450 (.A1(n_825), .A2(n_819), .ZN(n_606));
   NOR2_X1 i_451 (.A1(n_825), .A2(n_818), .ZN(n_607));
   NOR2_X1 i_452 (.A1(n_825), .A2(n_817), .ZN(n_608));
   NOR2_X1 i_453 (.A1(n_825), .A2(n_816), .ZN(n_609));
   NOR2_X1 i_454 (.A1(n_825), .A2(n_815), .ZN(n_610));
   NOR2_X1 i_456 (.A1(n_825), .A2(n_813), .ZN(n_612));
   NOR2_X1 i_459 (.A1(n_825), .A2(n_810), .ZN(n_615));
   NOR2_X1 i_460 (.A1(n_825), .A2(n_809), .ZN(n_616));
   INV_X1 i_462 (.A(n_619), .ZN(n_618));
   NOR2_X1 i_463 (.A1(n_824), .A2(n_820), .ZN(n_619));
   NOR2_X1 i_464 (.A1(n_824), .A2(n_819), .ZN(n_620));
   NOR2_X1 i_465 (.A1(n_824), .A2(n_818), .ZN(n_621));
   NOR2_X1 i_466 (.A1(n_824), .A2(n_817), .ZN(n_622));
   NOR2_X1 i_467 (.A1(n_824), .A2(n_816), .ZN(n_623));
   NOR2_X1 i_469 (.A1(n_824), .A2(n_814), .ZN(n_625));
   NOR2_X1 i_472 (.A1(n_824), .A2(n_811), .ZN(n_628));
   NOR2_X1 i_473 (.A1(n_824), .A2(n_810), .ZN(n_629));
   NOR2_X1 i_474 (.A1(n_823), .A2(n_821), .ZN(n_630));
   NOR2_X1 i_475 (.A1(n_823), .A2(n_820), .ZN(n_631));
   NOR2_X1 i_476 (.A1(n_823), .A2(n_819), .ZN(n_632));
   NOR2_X1 i_477 (.A1(n_823), .A2(n_818), .ZN(n_633));
   NOR2_X1 i_478 (.A1(n_823), .A2(n_817), .ZN(n_634));
   NOR2_X1 i_480 (.A1(n_823), .A2(n_815), .ZN(n_636));
   NOR2_X1 i_481 (.A1(n_823), .A2(n_814), .ZN(n_637));
   NOR2_X1 i_483 (.A1(n_823), .A2(n_812), .ZN(n_639));
   INV_X1 i_485 (.A(n_641), .ZN(mult[1]));
   OAI21_X1 i_486 (.A(n_780), .B1(n_783), .B2(n_782), .ZN(n_641));
   XOR2_X1 i_487 (.A(n_780), .B(n_642), .Z(mult[2]));
   OAI21_X1 i_488 (.A(n_779), .B1(n_0), .B2(n_785), .ZN(n_642));
   XNOR2_X1 i_489 (.A(n_778), .B(n_643), .ZN(mult[3]));
   OAI21_X1 i_490 (.A(n_786), .B1(n_2), .B2(n_4), .ZN(n_643));
   XOR2_X1 i_491 (.A(n_776), .B(n_644), .Z(mult[4]));
   XOR2_X1 i_492 (.A(n_6), .B(n_10), .Z(n_644));
   XOR2_X1 i_493 (.A(n_775), .B(n_651), .Z(mult[5]));
   XOR2_X1 i_494 (.A(n_650), .B(n_647), .Z(mult[6]));
   XOR2_X1 i_495 (.A(n_648), .B(n_645), .Z(mult[7]));
   NOR2_X1 i_496 (.A1(n_772), .A2(n_763), .ZN(n_645));
   XNOR2_X1 i_497 (.A(n_652), .B(n_646), .ZN(mult[8]));
   OAI22_X1 i_498 (.A1(n_38), .A2(n_40), .B1(n_763), .B2(n_648), .ZN(n_646));
   AOI21_X1 i_499 (.A(n_773), .B1(n_26), .B2(n_28), .ZN(n_647));
   AOI21_X1 i_500 (.A(n_773), .B1(n_767), .B2(n_649), .ZN(n_648));
   INV_X1 i_501 (.A(n_650), .ZN(n_649));
   AOI21_X1 i_502 (.A(n_770), .B1(n_775), .B2(n_768), .ZN(n_650));
   OAI21_X1 i_503 (.A(n_768), .B1(n_16), .B2(n_18), .ZN(n_651));
   NOR2_X1 i_504 (.A1(n_774), .A2(n_765), .ZN(n_652));
   XOR2_X1 i_505 (.A(n_761), .B(n_659), .Z(mult[9]));
   XOR2_X1 i_506 (.A(n_658), .B(n_655), .Z(mult[10]));
   XOR2_X1 i_507 (.A(n_656), .B(n_653), .Z(mult[11]));
   NOR2_X1 i_508 (.A1(n_758), .A2(n_749), .ZN(n_653));
   XNOR2_X1 i_509 (.A(n_660), .B(n_654), .ZN(mult[12]));
   OAI22_X1 i_510 (.A1(n_106), .A2(n_108), .B1(n_749), .B2(n_656), .ZN(n_654));
   AOI21_X1 i_511 (.A(n_759), .B1(n_86), .B2(n_88), .ZN(n_655));
   AOI21_X1 i_512 (.A(n_759), .B1(n_753), .B2(n_657), .ZN(n_656));
   INV_X1 i_513 (.A(n_658), .ZN(n_657));
   AOI21_X1 i_514 (.A(n_756), .B1(n_761), .B2(n_754), .ZN(n_658));
   OAI21_X1 i_515 (.A(n_754), .B1(n_68), .B2(n_70), .ZN(n_659));
   NOR2_X1 i_516 (.A1(n_760), .A2(n_751), .ZN(n_660));
   XOR2_X1 i_517 (.A(n_747), .B(n_667), .Z(mult[13]));
   XOR2_X1 i_518 (.A(n_666), .B(n_663), .Z(mult[14]));
   XOR2_X1 i_519 (.A(n_664), .B(n_661), .Z(mult[15]));
   NOR2_X1 i_520 (.A1(n_744), .A2(n_735), .ZN(n_661));
   XNOR2_X1 i_521 (.A(n_668), .B(n_662), .ZN(mult[16]));
   OAI22_X1 i_522 (.A1(n_177), .A2(n_198), .B1(n_735), .B2(n_664), .ZN(n_662));
   AOI21_X1 i_523 (.A(n_745), .B1(n_174), .B2(n_176), .ZN(n_663));
   AOI21_X1 i_524 (.A(n_745), .B1(n_739), .B2(n_665), .ZN(n_664));
   INV_X1 i_525 (.A(n_666), .ZN(n_665));
   AOI21_X1 i_526 (.A(n_742), .B1(n_747), .B2(n_740), .ZN(n_666));
   OAI21_X1 i_527 (.A(n_740), .B1(n_152), .B2(n_154), .ZN(n_667));
   NOR2_X1 i_528 (.A1(n_746), .A2(n_737), .ZN(n_668));
   XOR2_X1 i_529 (.A(n_733), .B(n_675), .Z(mult[17]));
   XOR2_X1 i_530 (.A(n_674), .B(n_671), .Z(mult[18]));
   XOR2_X1 i_531 (.A(n_672), .B(n_669), .Z(mult[19]));
   NOR2_X1 i_532 (.A1(n_730), .A2(n_721), .ZN(n_669));
   XNOR2_X1 i_533 (.A(n_676), .B(n_670), .ZN(mult[20]));
   OAI22_X1 i_534 (.A1(n_253), .A2(n_266), .B1(n_721), .B2(n_672), .ZN(n_670));
   AOI21_X1 i_535 (.A(n_731), .B1(n_237), .B2(n_252), .ZN(n_671));
   AOI21_X1 i_536 (.A(n_731), .B1(n_725), .B2(n_673), .ZN(n_672));
   INV_X1 i_537 (.A(n_674), .ZN(n_673));
   AOI21_X1 i_538 (.A(n_728), .B1(n_733), .B2(n_726), .ZN(n_674));
   OAI21_X1 i_539 (.A(n_726), .B1(n_219), .B2(n_236), .ZN(n_675));
   NOR2_X1 i_540 (.A1(n_732), .A2(n_723), .ZN(n_676));
   XOR2_X1 i_541 (.A(n_719), .B(n_683), .Z(mult[21]));
   XOR2_X1 i_542 (.A(n_682), .B(n_679), .Z(mult[22]));
   XOR2_X1 i_543 (.A(n_680), .B(n_677), .Z(mult[23]));
   NOR2_X1 i_544 (.A1(n_716), .A2(n_707), .ZN(n_677));
   XNOR2_X1 i_545 (.A(n_684), .B(n_678), .ZN(mult[24]));
   OAI22_X1 i_546 (.A1(n_297), .A2(n_302), .B1(n_707), .B2(n_680), .ZN(n_678));
   AOI21_X1 i_547 (.A(n_717), .B1(n_289), .B2(n_296), .ZN(n_679));
   AOI21_X1 i_548 (.A(n_717), .B1(n_711), .B2(n_681), .ZN(n_680));
   INV_X1 i_549 (.A(n_682), .ZN(n_681));
   AOI21_X1 i_550 (.A(n_714), .B1(n_719), .B2(n_712), .ZN(n_682));
   OAI21_X1 i_551 (.A(n_712), .B1(n_279), .B2(n_288), .ZN(n_683));
   NOR2_X1 i_552 (.A1(n_718), .A2(n_709), .ZN(n_684));
   XOR2_X1 i_553 (.A(n_705), .B(n_693), .Z(mult[25]));
   AOI22_X1 i_554 (.A1(n_692), .A2(n_689), .B1(n_691), .B2(n_690), .ZN(mult[26]));
   NOR2_X1 i_562 (.A1(n_792), .A2(n_700), .ZN(n_690));
   OR2_X1 i_565 (.A1(n_704), .A2(n_701), .ZN(n_693));
   INV_X1 i_567 (.A(n_695), .ZN(mult[29]));
   AOI21_X1 i_568 (.A(n_793), .B1(n_702), .B2(n_696), .ZN(n_695));
   AOI211_X1 i_569 (.A(n_698), .B(n_697), .C1(n_788), .C2(n_699), .ZN(n_696));
   AND2_X1 i_571 (.A1(n_805), .A2(n_794), .ZN(n_698));
   OR2_X1 i_572 (.A1(n_701), .A2(n_700), .ZN(n_699));
   NAND2_X1 i_575 (.A1(n_788), .A2(n_703), .ZN(n_702));
   INV_X1 i_580 (.A(n_708), .ZN(n_707));
   NAND2_X1 i_581 (.A1(n_297), .A2(n_302), .ZN(n_708));
   NAND2_X1 i_584 (.A1(n_289), .A2(n_296), .ZN(n_711));
   NAND2_X1 i_585 (.A1(n_279), .A2(n_288), .ZN(n_712));
   NOR2_X1 i_589 (.A1(n_297), .A2(n_302), .ZN(n_716));
   NOR2_X1 i_590 (.A1(n_289), .A2(n_296), .ZN(n_717));
   NOR2_X1 i_591 (.A1(n_303), .A2(n_306), .ZN(n_718));
   INV_X1 i_594 (.A(n_722), .ZN(n_721));
   NAND2_X1 i_595 (.A1(n_253), .A2(n_266), .ZN(n_722));
   NAND2_X1 i_598 (.A1(n_237), .A2(n_252), .ZN(n_725));
   NAND2_X1 i_599 (.A1(n_219), .A2(n_236), .ZN(n_726));
   NOR2_X1 i_603 (.A1(n_253), .A2(n_266), .ZN(n_730));
   NOR2_X1 i_604 (.A1(n_237), .A2(n_252), .ZN(n_731));
   NOR2_X1 i_605 (.A1(n_267), .A2(n_278), .ZN(n_732));
   INV_X1 i_608 (.A(n_736), .ZN(n_735));
   NAND2_X1 i_609 (.A1(n_177), .A2(n_198), .ZN(n_736));
   INV_X1 i_622 (.A(n_750), .ZN(n_749));
   INV_X1 i_636 (.A(n_764), .ZN(n_763));
   NAND2_X1 i_649 (.A1(n_786), .A2(n_777), .ZN(n_776));
   OAI21_X1 i_650 (.A(n_778), .B1(n_2), .B2(n_4), .ZN(n_777));
   AOI21_X1 i_651 (.A(n_784), .B1(n_780), .B2(n_779), .ZN(n_778));
   NAND2_X1 i_652 (.A1(n_0), .A2(n_785), .ZN(n_779));
   NAND2_X1 i_653 (.A1(mult[0]), .A2(n_781), .ZN(n_780));
   NOR2_X1 i_655 (.A1(n_823), .A2(n_808), .ZN(mult[0]));
   NOR2_X1 i_656 (.A1(n_823), .A2(n_809), .ZN(n_782));
   NOR2_X1 i_657 (.A1(n_824), .A2(n_808), .ZN(n_783));
   NOR2_X1 i_658 (.A1(n_0), .A2(n_785), .ZN(n_784));
   NOR2_X1 i_659 (.A1(n_823), .A2(n_810), .ZN(n_785));
   NAND2_X1 i_660 (.A1(n_2), .A2(n_4), .ZN(n_786));
   AND2_X1 i_661 (.A1(n_6), .A2(n_10), .ZN(n_787));
   AND2_X1 i_663 (.A1(n_806), .A2(n_790), .ZN(n_789));
   XOR2_X1 i_664 (.A(n_795), .B(n_791), .Z(n_790));
   NOR2_X1 i_665 (.A1(n_803), .A2(n_800), .ZN(n_791));
   NOR2_X1 i_666 (.A1(n_309), .A2(n_310), .ZN(n_792));
   NOR2_X1 i_667 (.A1(n_805), .A2(n_794), .ZN(n_793));
   OAI21_X1 i_668 (.A(n_804), .B1(n_800), .B2(n_795), .ZN(n_794));
   AOI21_X1 i_669 (.A(n_799), .B1(n_797), .B2(n_796), .ZN(n_795));
   NAND2_X1 i_670 (.A1(operand2[14]), .A2(operand1[12]), .ZN(n_796));
   INV_X1 i_671 (.A(n_798), .ZN(n_797));
   NOR3_X1 i_672 (.A1(n_835), .A2(n_822), .A3(n_802), .ZN(n_798));
   AOI21_X1 i_673 (.A(n_801), .B1(operand2[12]), .B2(operand1[14]), .ZN(n_799));
   NOR3_X1 i_674 (.A1(n_837), .A2(n_822), .A3(n_801), .ZN(n_800));
   INV_X1 i_675 (.A(n_802), .ZN(n_801));
   NOR2_X1 i_676 (.A1(n_836), .A2(n_821), .ZN(n_802));
   INV_X1 i_677 (.A(n_804), .ZN(n_803));
   OAI22_X1 i_678 (.A1(n_837), .A2(n_821), .B1(n_836), .B2(n_822), .ZN(n_804));
   NOR2_X1 i_679 (.A1(n_837), .A2(n_822), .ZN(n_805));
   INV_X1 i_680 (.A(n_311), .ZN(n_806));
   INV_X1 i_681 (.A(n_183), .ZN(n_807));
   INV_X1 i_691 (.A(operand1[9]), .ZN(n_817));
   INV_X1 i_692 (.A(operand1[10]), .ZN(n_818));
   INV_X1 i_693 (.A(operand1[11]), .ZN(n_819));
   INV_X1 i_694 (.A(operand1[12]), .ZN(n_820));
   INV_X1 i_695 (.A(operand1[13]), .ZN(n_821));
   INV_X1 i_696 (.A(operand1[14]), .ZN(n_822));
   INV_X1 i_703 (.A(operand2[6]), .ZN(n_829));
   INV_X1 i_704 (.A(operand2[7]), .ZN(n_830));
   INV_X1 i_705 (.A(operand2[8]), .ZN(n_831));
   INV_X1 i_706 (.A(operand2[9]), .ZN(n_832));
   INV_X1 i_707 (.A(operand2[10]), .ZN(n_833));
   INV_X1 i_708 (.A(operand2[11]), .ZN(n_834));
   INV_X1 i_709 (.A(operand2[12]), .ZN(n_835));
   INV_X1 i_710 (.A(operand2[13]), .ZN(n_836));
   INV_X1 i_711 (.A(operand2[14]), .ZN(n_837));
   NAND2_X1 i_420 (.A1(n_106), .A2(n_108), .ZN(n_750));
   INV_X1 i_423 (.A(n_852), .ZN(n_701));
   INV_X1 i_432 (.A(n_839), .ZN(n_703));
   NOR2_X1 i_435 (.A1(n_789), .A2(n_792), .ZN(n_788));
   INV_X1 i_444 (.A(n_690), .ZN(n_689));
   INV_X1 i_446 (.A(n_691), .ZN(n_692));
   INV_X1 i_447 (.A(n_854), .ZN(n_709));
   NOR2_X1 i_455 (.A1(n_279), .A2(n_288), .ZN(n_714));
   INV_X1 i_457 (.A(n_860), .ZN(n_719));
   INV_X1 i_458 (.A(n_863), .ZN(n_723));
   INV_X1 i_461 (.A(n_872), .ZN(n_733));
   INV_X1 i_468 (.A(n_875), .ZN(n_746));
   INV_X1 i_470 (.A(n_902), .ZN(n_742));
   INV_X1 i_471 (.A(n_910), .ZN(n_745));
   NOR2_X1 i_479 (.A1(n_177), .A2(n_198), .ZN(n_744));
   INV_X1 i_482 (.A(n_882), .ZN(n_747));
   INV_X1 i_484 (.A(n_883), .ZN(n_751));
   INV_X1 i_555 (.A(n_899), .ZN(n_760));
   NOR2_X1 i_556 (.A1(n_70), .A2(n_68), .ZN(n_756));
   INV_X1 i_557 (.A(n_890), .ZN(n_761));
   INV_X1 i_558 (.A(n_892), .ZN(n_765));
   INV_X1 i_559 (.A(operand2[5]), .ZN(n_828));
   INV_X1 i_560 (.A(operand1[0]), .ZN(n_808));
   INV_X1 i_561 (.A(operand1[2]), .ZN(n_810));
   INV_X1 i_563 (.A(operand2[2]), .ZN(n_825));
   INV_X1 i_564 (.A(operand2[0]), .ZN(n_823));
   INV_X1 i_566 (.A(operand1[1]), .ZN(n_809));
   INV_X1 i_570 (.A(operand2[1]), .ZN(n_824));
   INV_X1 i_573 (.A(operand1[3]), .ZN(n_811));
   INV_X1 i_574 (.A(operand1[4]), .ZN(n_812));
   INV_X1 i_576 (.A(operand2[3]), .ZN(n_826));
   INV_X1 i_577 (.A(operand1[5]), .ZN(n_813));
   INV_X1 i_578 (.A(operand2[4]), .ZN(n_827));
   INV_X1 i_579 (.A(operand1[6]), .ZN(n_814));
   INV_X1 i_582 (.A(operand1[7]), .ZN(n_815));
   INV_X1 i_583 (.A(operand1[8]), .ZN(n_816));
   INV_X1 i_586 (.A(n_685), .ZN(n_635));
   NAND2_X1 i_587 (.A1(operand1[8]), .A2(operand2[0]), .ZN(n_685));
   INV_X1 i_588 (.A(n_686), .ZN(n_624));
   NAND2_X1 i_592 (.A1(operand2[1]), .A2(operand1[7]), .ZN(n_686));
   INV_X1 i_593 (.A(n_687), .ZN(n_611));
   NAND2_X1 i_596 (.A1(operand2[2]), .A2(operand1[6]), .ZN(n_687));
   INV_X1 i_597 (.A(n_688), .ZN(n_600));
   NAND2_X1 i_600 (.A1(operand1[5]), .A2(operand2[3]), .ZN(n_688));
   INV_X1 i_601 (.A(n_694), .ZN(n_588));
   NAND2_X1 i_602 (.A1(operand2[4]), .A2(operand1[4]), .ZN(n_694));
   INV_X1 i_606 (.A(n_706), .ZN(n_576));
   NAND2_X1 i_607 (.A1(operand1[3]), .A2(operand2[5]), .ZN(n_706));
   INV_X1 i_610 (.A(n_710), .ZN(n_626));
   NAND2_X1 i_611 (.A1(operand2[1]), .A2(operand1[5]), .ZN(n_710));
   INV_X1 i_612 (.A(n_713), .ZN(n_613));
   NAND2_X1 i_613 (.A1(operand2[2]), .A2(operand1[4]), .ZN(n_713));
   INV_X1 i_614 (.A(n_715), .ZN(n_602));
   NAND2_X1 i_615 (.A1(operand1[3]), .A2(operand2[3]), .ZN(n_715));
   INV_X1 i_616 (.A(n_720), .ZN(n_638));
   NAND2_X1 i_617 (.A1(operand1[5]), .A2(operand2[0]), .ZN(n_720));
   INV_X1 i_618 (.A(n_724), .ZN(n_627));
   NAND2_X1 i_619 (.A1(operand2[1]), .A2(operand1[4]), .ZN(n_724));
   INV_X1 i_620 (.A(n_727), .ZN(n_614));
   NAND2_X1 i_621 (.A1(operand2[2]), .A2(operand1[3]), .ZN(n_727));
   INV_X1 i_623 (.A(n_729), .ZN(n_603));
   NAND2_X1 i_624 (.A1(operand1[2]), .A2(operand2[3]), .ZN(n_729));
   INV_X1 i_625 (.A(n_734), .ZN(n_591));
   NAND2_X1 i_626 (.A1(operand1[1]), .A2(operand2[4]), .ZN(n_734));
   INV_X1 i_627 (.A(n_738), .ZN(n_579));
   NAND2_X1 i_628 (.A1(operand1[0]), .A2(operand2[5]), .ZN(n_738));
   INV_X1 i_629 (.A(n_741), .ZN(n_640));
   NAND2_X1 i_630 (.A1(operand1[3]), .A2(operand2[0]), .ZN(n_741));
   INV_X1 i_631 (.A(n_743), .ZN(n_781));
   NAND2_X1 i_632 (.A1(operand2[1]), .A2(operand1[1]), .ZN(n_743));
   INV_X1 i_633 (.A(n_748), .ZN(n_617));
   NAND2_X1 i_634 (.A1(operand2[2]), .A2(operand1[0]), .ZN(n_748));
   INV_X1 i_635 (.A(n_752), .ZN(mult[27]));
   NAND2_X1 i_637 (.A1(n_769), .A2(n_755), .ZN(n_752));
   NAND3_X1 i_638 (.A1(n_757), .A2(n_766), .A3(n_844), .ZN(n_755));
   NAND2_X1 i_639 (.A1(n_691), .A2(n_762), .ZN(n_757));
   INV_X1 i_640 (.A(n_838), .ZN(n_762));
   INV_X1 i_641 (.A(n_845), .ZN(n_766));
   OAI21_X1 i_642 (.A(n_845), .B1(n_771), .B2(n_700), .ZN(n_769));
   AOI21_X1 i_643 (.A(n_838), .B1(n_839), .B2(n_852), .ZN(n_771));
   NOR2_X1 i_644 (.A1(n_309), .A2(n_310), .ZN(n_838));
   OAI21_X1 i_645 (.A(n_840), .B1(n_841), .B2(n_853), .ZN(n_839));
   INV_X1 i_646 (.A(n_704), .ZN(n_840));
   AOI21_X1 i_647 (.A(n_858), .B1(n_842), .B2(n_866), .ZN(n_841));
   AOI21_X1 i_648 (.A(n_862), .B1(n_843), .B2(n_865), .ZN(n_842));
   NOR2_X1 i_654 (.A1(n_731), .A2(n_869), .ZN(n_843));
   INV_X1 i_662 (.A(n_844), .ZN(n_700));
   NAND2_X1 i_682 (.A1(n_309), .A2(n_310), .ZN(n_844));
   NOR2_X1 i_683 (.A1(n_789), .A2(n_697), .ZN(n_845));
   NAND2_X1 i_684 (.A1(n_846), .A2(n_848), .ZN(mult[28]));
   NAND2_X1 i_685 (.A1(n_847), .A2(n_915), .ZN(n_846));
   OAI21_X1 i_686 (.A(n_849), .B1(n_691), .B2(n_850), .ZN(n_847));
   OAI211_X1 i_687 (.A(n_914), .B(n_849), .C1(n_691), .C2(n_850), .ZN(n_848));
   OAI21_X1 i_688 (.A(n_851), .B1(n_789), .B2(n_792), .ZN(n_849));
   NAND2_X1 i_689 (.A1(n_690), .A2(n_851), .ZN(n_850));
   INV_X1 i_690 (.A(n_697), .ZN(n_851));
   NOR2_X1 i_697 (.A1(n_806), .A2(n_790), .ZN(n_697));
   OAI21_X1 i_698 (.A(n_852), .B1(n_705), .B2(n_704), .ZN(n_691));
   NAND2_X1 i_699 (.A1(n_307), .A2(n_308), .ZN(n_852));
   NOR2_X1 i_700 (.A1(n_307), .A2(n_308), .ZN(n_704));
   AOI21_X1 i_701 (.A(n_853), .B1(n_860), .B2(n_857), .ZN(n_705));
   OAI211_X1 i_702 (.A(n_855), .B(n_854), .C1(n_718), .C2(n_708), .ZN(n_853));
   NAND2_X1 i_712 (.A1(n_303), .A2(n_306), .ZN(n_854));
   NAND2_X1 i_713 (.A1(n_859), .A2(n_856), .ZN(n_855));
   NAND2_X1 i_714 (.A1(n_712), .A2(n_711), .ZN(n_856));
   INV_X1 i_715 (.A(n_858), .ZN(n_857));
   OAI21_X1 i_716 (.A(n_859), .B1(n_279), .B2(n_288), .ZN(n_858));
   NOR3_X1 i_717 (.A1(n_717), .A2(n_716), .A3(n_718), .ZN(n_859));
   NAND3_X1 i_718 (.A1(n_866), .A2(n_864), .A3(n_861), .ZN(n_860));
   INV_X1 i_719 (.A(n_862), .ZN(n_861));
   OAI21_X1 i_720 (.A(n_863), .B1(n_722), .B2(n_732), .ZN(n_862));
   NAND2_X1 i_721 (.A1(n_267), .A2(n_278), .ZN(n_863));
   NAND3_X1 i_722 (.A1(n_913), .A2(n_868), .A3(n_865), .ZN(n_864));
   NAND2_X1 i_723 (.A1(n_725), .A2(n_726), .ZN(n_865));
   NAND4_X1 i_724 (.A1(n_872), .A2(n_913), .A3(n_868), .A4(n_867), .ZN(n_866));
   INV_X1 i_725 (.A(n_728), .ZN(n_867));
   NOR2_X1 i_726 (.A1(n_236), .A2(n_219), .ZN(n_728));
   INV_X1 i_727 (.A(n_869), .ZN(n_868));
   NAND2_X1 i_728 (.A1(n_871), .A2(n_870), .ZN(n_869));
   INV_X1 i_729 (.A(n_732), .ZN(n_870));
   INV_X1 i_730 (.A(n_730), .ZN(n_871));
   NAND3_X1 i_731 (.A1(n_877), .A2(n_879), .A3(n_873), .ZN(n_872));
   AOI21_X1 i_732 (.A(n_737), .B1(n_876), .B2(n_875), .ZN(n_873));
   INV_X1 i_733 (.A(n_874), .ZN(n_737));
   NAND2_X1 i_734 (.A1(n_218), .A2(n_199), .ZN(n_874));
   NAND2_X1 i_735 (.A1(n_906), .A2(n_908), .ZN(n_875));
   INV_X1 i_736 (.A(n_736), .ZN(n_876));
   NAND3_X1 i_737 (.A1(n_878), .A2(n_905), .A3(n_910), .ZN(n_877));
   NAND2_X1 i_738 (.A1(n_739), .A2(n_740), .ZN(n_878));
   NAND2_X1 i_739 (.A1(n_176), .A2(n_174), .ZN(n_739));
   NAND2_X1 i_740 (.A1(n_154), .A2(n_152), .ZN(n_740));
   NAND3_X1 i_741 (.A1(n_905), .A2(n_910), .A3(n_880), .ZN(n_879));
   INV_X1 i_742 (.A(n_881), .ZN(n_880));
   NAND2_X1 i_743 (.A1(n_882), .A2(n_902), .ZN(n_881));
   NAND4_X1 i_744 (.A1(n_887), .A2(n_885), .A3(n_884), .A4(n_883), .ZN(n_882));
   NAND2_X1 i_745 (.A1(n_130), .A2(n_128), .ZN(n_883));
   NAND3_X1 i_746 (.A1(n_899), .A2(n_106), .A3(n_108), .ZN(n_884));
   NAND3_X1 i_747 (.A1(n_898), .A2(n_899), .A3(n_886), .ZN(n_885));
   NAND2_X1 i_748 (.A1(n_753), .A2(n_754), .ZN(n_886));
   NAND2_X1 i_749 (.A1(n_88), .A2(n_86), .ZN(n_753));
   NAND2_X1 i_750 (.A1(n_70), .A2(n_68), .ZN(n_754));
   NAND3_X1 i_751 (.A1(n_898), .A2(n_899), .A3(n_888), .ZN(n_887));
   INV_X1 i_752 (.A(n_889), .ZN(n_888));
   OAI21_X1 i_753 (.A(n_890), .B1(n_68), .B2(n_70), .ZN(n_889));
   NAND4_X1 i_754 (.A1(n_891), .A2(n_895), .A3(n_893), .A4(n_892), .ZN(n_890));
   OR2_X1 i_755 (.A1(n_774), .A2(n_764), .ZN(n_891));
   NAND2_X1 i_756 (.A1(n_38), .A2(n_40), .ZN(n_764));
   NOR2_X1 i_757 (.A1(n_54), .A2(n_52), .ZN(n_774));
   NAND2_X1 i_758 (.A1(n_54), .A2(n_52), .ZN(n_892));
   OAI211_X1 i_759 (.A(n_897), .B(n_894), .C1(n_52), .C2(n_54), .ZN(n_893));
   NAND2_X1 i_760 (.A1(n_767), .A2(n_768), .ZN(n_894));
   NAND2_X1 i_761 (.A1(n_28), .A2(n_26), .ZN(n_767));
   NAND2_X1 i_762 (.A1(n_18), .A2(n_16), .ZN(n_768));
   OAI211_X1 i_763 (.A(n_897), .B(n_896), .C1(n_52), .C2(n_54), .ZN(n_895));
   NOR2_X1 i_764 (.A1(n_775), .A2(n_770), .ZN(n_896));
   NOR2_X1 i_765 (.A1(n_18), .A2(n_16), .ZN(n_770));
   OAI22_X1 i_766 (.A1(n_787), .A2(n_776), .B1(n_6), .B2(n_10), .ZN(n_775));
   NOR2_X1 i_767 (.A1(n_772), .A2(n_773), .ZN(n_897));
   NOR2_X1 i_768 (.A1(n_38), .A2(n_40), .ZN(n_772));
   NOR2_X1 i_769 (.A1(n_28), .A2(n_26), .ZN(n_773));
   NOR2_X1 i_770 (.A1(n_758), .A2(n_759), .ZN(n_898));
   NOR2_X1 i_771 (.A1(n_88), .A2(n_86), .ZN(n_759));
   NOR2_X1 i_772 (.A1(n_106), .A2(n_108), .ZN(n_758));
   NAND2_X1 i_773 (.A1(n_900), .A2(n_901), .ZN(n_899));
   INV_X1 i_774 (.A(n_130), .ZN(n_900));
   INV_X1 i_775 (.A(n_128), .ZN(n_901));
   NAND2_X1 i_776 (.A1(n_903), .A2(n_904), .ZN(n_902));
   INV_X1 i_777 (.A(n_154), .ZN(n_903));
   INV_X1 i_778 (.A(n_152), .ZN(n_904));
   AOI22_X1 i_779 (.A1(n_908), .A2(n_906), .B1(n_909), .B2(n_907), .ZN(n_905));
   INV_X1 i_780 (.A(n_218), .ZN(n_906));
   INV_X1 i_781 (.A(n_198), .ZN(n_907));
   INV_X1 i_782 (.A(n_199), .ZN(n_908));
   INV_X1 i_783 (.A(n_177), .ZN(n_909));
   NAND2_X1 i_784 (.A1(n_911), .A2(n_912), .ZN(n_910));
   INV_X1 i_785 (.A(n_176), .ZN(n_911));
   INV_X1 i_786 (.A(n_174), .ZN(n_912));
   INV_X1 i_787 (.A(n_731), .ZN(n_913));
   INV_X1 i_788 (.A(n_915), .ZN(n_914));
   NOR2_X1 i_789 (.A1(n_698), .A2(n_793), .ZN(n_915));
endmodule

module second_stage(operand1, operand2, clk, enable, negative_product, 
      next_stage_enable, negative_product_third_stage, product);
   input [14:0]operand1;
   input [14:0]operand2;
   input clk;
   input enable;
   input negative_product;
   output next_stage_enable;
   output negative_product_third_stage;
   output [29:0]product;

   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_0;
   wire n_0_2;

   CLKGATETST_X1 clk_gate_product_reg (.CK(clk), .E(1'b1), .SE(1'b0), .GCK(n_0_1));
   DFF_X1 \product_reg[29]  (.D(n_0_0), .CK(n_0_1), .Q(product[29]), .QN());
   DFF_X1 \product_reg[28]  (.D(n_0_31), .CK(n_0_1), .Q(product[28]), .QN());
   DFF_X1 \product_reg[27]  (.D(n_0_30), .CK(n_0_1), .Q(product[27]), .QN());
   DFF_X1 \product_reg[26]  (.D(n_0_29), .CK(n_0_1), .Q(product[26]), .QN());
   DFF_X1 \product_reg[25]  (.D(n_0_28), .CK(n_0_1), .Q(product[25]), .QN());
   DFF_X1 \product_reg[24]  (.D(n_0_27), .CK(n_0_1), .Q(product[24]), .QN());
   DFF_X1 \product_reg[23]  (.D(n_0_26), .CK(n_0_1), .Q(product[23]), .QN());
   DFF_X1 \product_reg[22]  (.D(n_0_25), .CK(n_0_1), .Q(product[22]), .QN());
   DFF_X1 \product_reg[21]  (.D(n_0_24), .CK(n_0_1), .Q(product[21]), .QN());
   DFF_X1 \product_reg[20]  (.D(n_0_23), .CK(n_0_1), .Q(product[20]), .QN());
   DFF_X1 \product_reg[19]  (.D(n_0_22), .CK(n_0_1), .Q(product[19]), .QN());
   DFF_X1 \product_reg[18]  (.D(n_0_21), .CK(n_0_1), .Q(product[18]), .QN());
   DFF_X1 \product_reg[17]  (.D(n_0_20), .CK(n_0_1), .Q(product[17]), .QN());
   DFF_X1 \product_reg[16]  (.D(n_0_19), .CK(n_0_1), .Q(product[16]), .QN());
   DFF_X1 \product_reg[15]  (.D(n_0_18), .CK(n_0_1), .Q(product[15]), .QN());
   DFF_X1 \product_reg[14]  (.D(n_0_17), .CK(n_0_1), .Q(product[14]), .QN());
   DFF_X1 \product_reg[13]  (.D(n_0_16), .CK(n_0_1), .Q(product[13]), .QN());
   DFF_X1 \product_reg[12]  (.D(n_0_15), .CK(n_0_1), .Q(product[12]), .QN());
   DFF_X1 \product_reg[11]  (.D(n_0_14), .CK(n_0_1), .Q(product[11]), .QN());
   DFF_X1 \product_reg[10]  (.D(n_0_13), .CK(n_0_1), .Q(product[10]), .QN());
   DFF_X1 \product_reg[9]  (.D(n_0_12), .CK(n_0_1), .Q(product[9]), .QN());
   DFF_X1 \product_reg[8]  (.D(n_0_11), .CK(n_0_1), .Q(product[8]), .QN());
   DFF_X1 \product_reg[7]  (.D(n_0_10), .CK(n_0_1), .Q(product[7]), .QN());
   DFF_X1 \product_reg[6]  (.D(n_0_9), .CK(n_0_1), .Q(product[6]), .QN());
   DFF_X1 \product_reg[5]  (.D(n_0_8), .CK(n_0_1), .Q(product[5]), .QN());
   DFF_X1 \product_reg[4]  (.D(n_0_7), .CK(n_0_1), .Q(product[4]), .QN());
   DFF_X1 \product_reg[3]  (.D(n_0_6), .CK(n_0_1), .Q(product[3]), .QN());
   DFF_X1 \product_reg[2]  (.D(n_0_5), .CK(n_0_1), .Q(product[2]), .QN());
   DFF_X2 \product_reg[1]  (.D(n_0_4), .CK(n_0_1), .Q(product[1]), .QN());
   DFF_X2 \product_reg[0]  (.D(n_0_3), .CK(n_0_1), .Q(product[0]), .QN());
   DFF_X1 negative_product_third_stage_reg (.D(negative_product), .CK(n_0_2), 
      .Q(negative_product_third_stage), .QN());
   datapath__0_4 i_0_1 (.operand2(operand2), .operand1(operand1), .mult({n_0_0, 
      n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, 
      n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
      n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, 
      n_0_3}));
   INV_X1 i_0_0_0 (.A(clk), .ZN(n_0_2));
endmodule

module datapath__0_71(product, minus);
   input [29:0]product;
   output [29:0]minus;

   AOI21_X1 i_0 (.A(n_58), .B1(product[1]), .B2(product[0]), .ZN(minus[1]));
   AOI21_X1 i_1 (.A(n_56), .B1(product[2]), .B2(n_57), .ZN(minus[2]));
   AOI21_X1 i_2 (.A(n_54), .B1(product[3]), .B2(n_55), .ZN(minus[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(product[4]), .B2(n_53), .ZN(minus[4]));
   AOI21_X1 i_4 (.A(n_3), .B1(product[5]), .B2(n_4), .ZN(minus[5]));
   AOI21_X1 i_5 (.A(n_1), .B1(product[6]), .B2(n_2), .ZN(minus[6]));
   AOI21_X1 i_6 (.A(n_51), .B1(product[7]), .B2(n_0), .ZN(minus[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   NOR2_X1 i_8 (.A1(n_53), .A2(n_52), .ZN(n_1));
   INV_X1 i_9 (.A(n_3), .ZN(n_2));
   NOR2_X1 i_10 (.A1(product[5]), .A2(n_4), .ZN(n_3));
   INV_X1 i_11 (.A(n_5), .ZN(n_4));
   NOR2_X1 i_12 (.A1(product[4]), .A2(n_53), .ZN(n_5));
   AOI21_X1 i_13 (.A(n_11), .B1(product[8]), .B2(n_50), .ZN(minus[8]));
   AOI21_X1 i_14 (.A(n_9), .B1(product[9]), .B2(n_10), .ZN(minus[9]));
   AOI21_X1 i_15 (.A(n_7), .B1(product[10]), .B2(n_8), .ZN(minus[10]));
   AOI21_X1 i_16 (.A(n_48), .B1(product[11]), .B2(n_6), .ZN(minus[11]));
   INV_X1 i_17 (.A(n_7), .ZN(n_6));
   NOR2_X1 i_18 (.A1(n_50), .A2(n_49), .ZN(n_7));
   INV_X1 i_19 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_20 (.A1(product[9]), .A2(n_10), .ZN(n_9));
   INV_X1 i_21 (.A(n_11), .ZN(n_10));
   NOR2_X1 i_22 (.A1(product[8]), .A2(n_50), .ZN(n_11));
   AOI21_X1 i_23 (.A(n_17), .B1(product[12]), .B2(n_47), .ZN(minus[12]));
   AOI21_X1 i_24 (.A(n_15), .B1(product[13]), .B2(n_16), .ZN(minus[13]));
   AOI21_X1 i_25 (.A(n_13), .B1(product[14]), .B2(n_14), .ZN(minus[14]));
   AOI21_X1 i_26 (.A(n_45), .B1(product[15]), .B2(n_12), .ZN(minus[15]));
   INV_X1 i_27 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_28 (.A1(n_47), .A2(n_46), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   NOR2_X1 i_30 (.A1(product[13]), .A2(n_16), .ZN(n_15));
   INV_X1 i_31 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_32 (.A1(product[12]), .A2(n_47), .ZN(n_17));
   AOI21_X1 i_33 (.A(n_23), .B1(product[16]), .B2(n_44), .ZN(minus[16]));
   AOI21_X1 i_34 (.A(n_21), .B1(product[17]), .B2(n_22), .ZN(minus[17]));
   AOI21_X1 i_35 (.A(n_19), .B1(product[18]), .B2(n_20), .ZN(minus[18]));
   AOI21_X1 i_36 (.A(n_41), .B1(product[19]), .B2(n_18), .ZN(minus[19]));
   INV_X1 i_37 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_38 (.A1(n_44), .A2(n_42), .ZN(n_19));
   INV_X1 i_39 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_40 (.A1(product[17]), .A2(n_22), .ZN(n_21));
   INV_X1 i_41 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_42 (.A1(product[16]), .A2(n_44), .ZN(n_23));
   AOI21_X1 i_43 (.A(n_25), .B1(product[20]), .B2(n_40), .ZN(minus[20]));
   AOI21_X1 i_44 (.A(n_27), .B1(product[21]), .B2(n_24), .ZN(minus[21]));
   INV_X1 i_45 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_46 (.A1(product[20]), .A2(n_40), .ZN(n_25));
   AOI21_X1 i_47 (.A(n_39), .B1(product[22]), .B2(n_26), .ZN(minus[22]));
   INV_X1 i_48 (.A(n_27), .ZN(n_26));
   NOR3_X1 i_49 (.A1(product[21]), .A2(product[20]), .A3(n_40), .ZN(n_27));
   AOI21_X1 i_50 (.A(n_37), .B1(product[23]), .B2(n_38), .ZN(minus[23]));
   AOI21_X1 i_51 (.A(n_29), .B1(product[24]), .B2(n_36), .ZN(minus[24]));
   AOI21_X1 i_55 (.A(n_32), .B1(product[26]), .B2(n_30), .ZN(minus[26]));
   NOR2_X1 i_59 (.A1(n_43), .A2(n_36), .ZN(n_32));
   NAND2_X1 i_52 (.A1(n_29), .A2(n_33), .ZN(n_30));
   INV_X1 i_53 (.A(n_28), .ZN(n_29));
   XNOR2_X1 i_54 (.A(n_28), .B(n_33), .ZN(minus[25]));
   NAND2_X1 i_56 (.A1(n_37), .A2(n_31), .ZN(n_28));
   INV_X1 i_57 (.A(product[24]), .ZN(n_31));
   INV_X1 i_58 (.A(product[25]), .ZN(n_33));
   AOI21_X1 i_60 (.A(n_60), .B1(n_34), .B2(product[27]), .ZN(minus[27]));
   INV_X1 i_61 (.A(n_32), .ZN(n_34));
   XNOR2_X1 i_62 (.A(n_61), .B(n_79), .ZN(minus[28]));
   OR2_X1 i_69 (.A1(n_43), .A2(product[27]), .ZN(n_63));
   OR3_X1 i_70 (.A1(product[25]), .A2(product[24]), .A3(product[26]), .ZN(n_43));
   OR3_X1 i_76 (.A1(product[20]), .A2(product[21]), .A3(product[22]), .ZN(n_65));
   OR2_X1 i_80 (.A1(n_42), .A2(product[19]), .ZN(n_67));
   OR3_X1 i_81 (.A1(product[17]), .A2(product[16]), .A3(product[18]), .ZN(n_42));
   OR2_X1 i_85 (.A1(n_46), .A2(product[15]), .ZN(n_69));
   OR3_X1 i_86 (.A1(product[13]), .A2(product[12]), .A3(product[14]), .ZN(n_46));
   INV_X1 i_63 (.A(n_61), .ZN(n_60));
   NAND2_X1 i_64 (.A1(n_37), .A2(n_85), .ZN(n_61));
   INV_X1 i_65 (.A(n_40), .ZN(n_41));
   NAND2_X1 i_66 (.A1(n_45), .A2(n_82), .ZN(n_40));
   INV_X1 i_67 (.A(n_45), .ZN(n_44));
   INV_X1 i_68 (.A(n_50), .ZN(n_51));
   NAND2_X1 i_71 (.A1(n_73), .A2(n_54), .ZN(n_50));
   INV_X1 i_72 (.A(n_35), .ZN(minus[29]));
   NAND2_X1 i_73 (.A1(n_66), .A2(n_59), .ZN(n_35));
   NAND2_X1 i_74 (.A1(n_62), .A2(product[29]), .ZN(n_59));
   NAND4_X1 i_75 (.A1(n_39), .A2(n_79), .A3(n_84), .A4(n_85), .ZN(n_62));
   INV_X1 i_77 (.A(n_38), .ZN(n_39));
   NAND4_X1 i_78 (.A1(n_82), .A2(n_64), .A3(n_83), .A4(n_48), .ZN(n_38));
   INV_X1 i_79 (.A(n_47), .ZN(n_48));
   INV_X1 i_82 (.A(n_69), .ZN(n_64));
   NAND4_X1 i_83 (.A1(n_37), .A2(n_86), .A3(n_79), .A4(n_85), .ZN(n_66));
   INV_X1 i_84 (.A(n_36), .ZN(n_37));
   NAND4_X1 i_87 (.A1(n_45), .A2(n_84), .A3(n_83), .A4(n_82), .ZN(n_36));
   NOR2_X1 i_88 (.A1(n_69), .A2(n_47), .ZN(n_45));
   NAND3_X1 i_89 (.A1(n_73), .A2(n_68), .A3(n_54), .ZN(n_47));
   INV_X1 i_90 (.A(n_70), .ZN(n_68));
   OR2_X1 i_91 (.A1(n_49), .A2(product[11]), .ZN(n_70));
   NAND2_X1 i_92 (.A1(n_71), .A2(n_72), .ZN(n_49));
   NOR2_X1 i_93 (.A1(product[9]), .A2(product[10]), .ZN(n_71));
   INV_X1 i_94 (.A(product[8]), .ZN(n_72));
   INV_X1 i_95 (.A(n_74), .ZN(n_73));
   OR2_X1 i_96 (.A1(n_52), .A2(product[7]), .ZN(n_74));
   NAND2_X1 i_97 (.A1(n_75), .A2(n_76), .ZN(n_52));
   NOR2_X1 i_98 (.A1(product[5]), .A2(product[6]), .ZN(n_75));
   INV_X1 i_99 (.A(product[4]), .ZN(n_76));
   INV_X1 i_100 (.A(n_53), .ZN(n_54));
   NAND2_X1 i_101 (.A1(n_56), .A2(n_81), .ZN(n_53));
   INV_X1 i_102 (.A(n_55), .ZN(n_56));
   NAND2_X1 i_103 (.A1(n_58), .A2(n_80), .ZN(n_55));
   INV_X1 i_104 (.A(n_57), .ZN(n_58));
   NAND2_X1 i_105 (.A1(n_77), .A2(n_78), .ZN(n_57));
   INV_X1 i_106 (.A(product[0]), .ZN(n_77));
   INV_X1 i_107 (.A(product[1]), .ZN(n_78));
   INV_X1 i_108 (.A(product[2]), .ZN(n_80));
   INV_X1 i_109 (.A(product[3]), .ZN(n_81));
   INV_X1 i_110 (.A(n_67), .ZN(n_82));
   INV_X1 i_111 (.A(n_65), .ZN(n_83));
   INV_X1 i_112 (.A(product[23]), .ZN(n_84));
   INV_X1 i_113 (.A(n_63), .ZN(n_85));
   INV_X1 i_114 (.A(product[28]), .ZN(n_79));
   INV_X1 i_115 (.A(product[29]), .ZN(n_86));
endmodule

module third_stage(clk, enable, negative_product, product, C);
   input clk;
   input enable;
   input negative_product;
   input [29:0]product;
   output [30:0]C;

   datapath__0_71 i_1 (.product(product), .minus({n_28, n_27, n_26, n_25, n_24, 
      n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
      n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_0}));
   MUX2_X1 i_0_0 (.A(product[1]), .B(n_0), .S(negative_product), .Z(n_29));
   MUX2_X1 i_0_1 (.A(product[2]), .B(n_1), .S(negative_product), .Z(n_30));
   MUX2_X1 i_0_2 (.A(product[3]), .B(n_2), .S(negative_product), .Z(n_31));
   MUX2_X1 i_0_3 (.A(product[4]), .B(n_3), .S(negative_product), .Z(n_32));
   MUX2_X1 i_0_4 (.A(product[5]), .B(n_4), .S(negative_product), .Z(n_33));
   MUX2_X1 i_0_5 (.A(product[6]), .B(n_5), .S(negative_product), .Z(n_34));
   MUX2_X1 i_0_6 (.A(product[7]), .B(n_6), .S(negative_product), .Z(n_35));
   MUX2_X1 i_0_7 (.A(product[8]), .B(n_7), .S(negative_product), .Z(n_36));
   MUX2_X1 i_0_8 (.A(product[9]), .B(n_8), .S(negative_product), .Z(n_37));
   MUX2_X1 i_0_9 (.A(product[10]), .B(n_9), .S(negative_product), .Z(n_38));
   MUX2_X1 i_0_10 (.A(product[11]), .B(n_10), .S(negative_product), .Z(n_39));
   MUX2_X1 i_0_11 (.A(product[12]), .B(n_11), .S(negative_product), .Z(n_40));
   MUX2_X1 i_0_12 (.A(product[13]), .B(n_12), .S(negative_product), .Z(n_41));
   MUX2_X1 i_0_13 (.A(product[14]), .B(n_13), .S(negative_product), .Z(n_42));
   MUX2_X1 i_0_14 (.A(product[15]), .B(n_14), .S(negative_product), .Z(n_43));
   MUX2_X1 i_0_15 (.A(product[16]), .B(n_15), .S(negative_product), .Z(n_44));
   MUX2_X1 i_0_16 (.A(product[17]), .B(n_16), .S(negative_product), .Z(n_45));
   MUX2_X1 i_0_17 (.A(product[18]), .B(n_17), .S(negative_product), .Z(n_46));
   MUX2_X1 i_0_18 (.A(product[19]), .B(n_18), .S(negative_product), .Z(n_47));
   MUX2_X1 i_0_19 (.A(product[20]), .B(n_19), .S(negative_product), .Z(n_48));
   MUX2_X1 i_0_20 (.A(product[21]), .B(n_20), .S(negative_product), .Z(n_49));
   MUX2_X1 i_0_21 (.A(product[22]), .B(n_21), .S(negative_product), .Z(n_50));
   MUX2_X1 i_0_22 (.A(product[23]), .B(n_22), .S(negative_product), .Z(n_51));
   MUX2_X1 i_0_23 (.A(product[24]), .B(n_23), .S(negative_product), .Z(n_52));
   MUX2_X1 i_0_24 (.A(product[25]), .B(n_24), .S(negative_product), .Z(n_53));
   MUX2_X1 i_0_25 (.A(product[26]), .B(n_25), .S(negative_product), .Z(n_54));
   MUX2_X1 i_0_26 (.A(product[27]), .B(n_26), .S(negative_product), .Z(n_55));
   MUX2_X1 i_0_27 (.A(product[28]), .B(n_27), .S(negative_product), .Z(n_56));
   MUX2_X1 i_0_28 (.A(product[29]), .B(n_28), .S(negative_product), .Z(n_57));
   INV_X1 i_0_29 (.A(clk), .ZN(n_58));
   DFF_X1 \C_reg[30]  (.D(negative_product), .CK(n_58), .Q(C[30]), .QN());
   DFF_X1 \C_reg[29]  (.D(n_57), .CK(n_58), .Q(C[29]), .QN());
   DFF_X1 \C_reg[28]  (.D(n_56), .CK(n_58), .Q(C[28]), .QN());
   DFF_X1 \C_reg[27]  (.D(n_55), .CK(n_58), .Q(C[27]), .QN());
   DFF_X1 \C_reg[26]  (.D(n_54), .CK(n_58), .Q(C[26]), .QN());
   DFF_X1 \C_reg[25]  (.D(n_53), .CK(n_58), .Q(C[25]), .QN());
   DFF_X1 \C_reg[24]  (.D(n_52), .CK(n_58), .Q(C[24]), .QN());
   DFF_X1 \C_reg[23]  (.D(n_51), .CK(n_58), .Q(C[23]), .QN());
   DFF_X1 \C_reg[22]  (.D(n_50), .CK(n_58), .Q(C[22]), .QN());
   DFF_X1 \C_reg[21]  (.D(n_49), .CK(n_58), .Q(C[21]), .QN());
   DFF_X1 \C_reg[20]  (.D(n_48), .CK(n_58), .Q(C[20]), .QN());
   DFF_X1 \C_reg[19]  (.D(n_47), .CK(n_58), .Q(C[19]), .QN());
   DFF_X1 \C_reg[18]  (.D(n_46), .CK(n_58), .Q(C[18]), .QN());
   DFF_X1 \C_reg[17]  (.D(n_45), .CK(n_58), .Q(C[17]), .QN());
   DFF_X1 \C_reg[16]  (.D(n_44), .CK(n_58), .Q(C[16]), .QN());
   DFF_X1 \C_reg[15]  (.D(n_43), .CK(n_58), .Q(C[15]), .QN());
   DFF_X1 \C_reg[14]  (.D(n_42), .CK(n_58), .Q(C[14]), .QN());
   DFF_X1 \C_reg[13]  (.D(n_41), .CK(n_58), .Q(C[13]), .QN());
   DFF_X1 \C_reg[12]  (.D(n_40), .CK(n_58), .Q(C[12]), .QN());
   DFF_X1 \C_reg[11]  (.D(n_39), .CK(n_58), .Q(C[11]), .QN());
   DFF_X1 \C_reg[10]  (.D(n_38), .CK(n_58), .Q(C[10]), .QN());
   DFF_X1 \C_reg[9]  (.D(n_37), .CK(n_58), .Q(C[9]), .QN());
   DFF_X1 \C_reg[8]  (.D(n_36), .CK(n_58), .Q(C[8]), .QN());
   DFF_X1 \C_reg[7]  (.D(n_35), .CK(n_58), .Q(C[7]), .QN());
   DFF_X1 \C_reg[6]  (.D(n_34), .CK(n_58), .Q(C[6]), .QN());
   DFF_X1 \C_reg[5]  (.D(n_33), .CK(n_58), .Q(C[5]), .QN());
   DFF_X1 \C_reg[4]  (.D(n_32), .CK(n_58), .Q(C[4]), .QN());
   DFF_X1 \C_reg[3]  (.D(n_31), .CK(n_58), .Q(C[3]), .QN());
   DFF_X1 \C_reg[2]  (.D(n_30), .CK(n_58), .Q(C[2]), .QN());
   DFF_X1 \C_reg[1]  (.D(n_29), .CK(n_58), .Q(C[1]), .QN());
   DFF_X1 \C_reg[0]  (.D(product[0]), .CK(n_58), .Q(C[0]), .QN());
endmodule

module pipelined_multiplier(A, B, clk, enable, C);
   input [15:0]A;
   input [15:0]B;
   input clk;
   input enable;
   output [30:0]C;

   wire [14:0]operand2;
   wire [14:0]operand1;
   wire negative_product_second_stage;
   wire [29:0]product;
   wire negative_product_third_stage;

   first_stage stage1 (.A(A), .B(B), .clk(clk), .enable(enable), 
      .negative_product_second_stage(negative_product_second_stage), 
      .next_stage_enable(), .operand1(operand1), .operand2(operand2));
   second_stage stage2 (.operand1(operand1), .operand2(operand2), .clk(clk), 
      .enable(), .negative_product(negative_product_second_stage), 
      .next_stage_enable(), .negative_product_third_stage(
      negative_product_third_stage), .product(product));
   third_stage stage3 (.clk(clk), .enable(), .negative_product(
      negative_product_third_stage), .product(product), .C(C));
endmodule
